`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
X92hFfkJFYFA0DNyC8rGa5S4bBAysNK3be3Aq1AI2jPyJXBpPxitBV/MlxV68cS7dunjMuyUVVTm
sFS8vqPaKQ==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NSquXs3p89GeQ3RkBK97ec+jzL/3jLE91bL5RxgYC2QNnsgtW9bDgLYt63iAvB9laJZLHrJnsumd
x8cKjY/uR09nIcO6h+Yc5HM3p8BYNQTwheeyLpF9wfAbuwu+OAM3JGDRd+/c6K3Jq+xWJvXEBoTJ
CW+mb4WNCAe5CcE9gdE=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nffxmj8+kDVElG/S83a+wtOhybK7y3bsZG/5mNoMwCFy+djZy4sbzpzzqHgEZJvOgsThiijbJMak
DW9OArJcrDp05IX768z09/z6BvtLq9ErH8Zx9j/kG2lzttaJyZskOtLll5nAuWHV0puT3Dm1Rpnb
foaFmA9QJWjenm42rHtDqwRwXXVnt0i+dxFPernAOuuAUvPK+PTmdQZFmqgUpCg0aBnTfHD7I7rI
Mm6C7TP9Eup8qggKjPnrESUP3HMknTcvAdfEhElfQ09JRxbYJqW3xOzik1K9Oz9VQxX9lPCkqe6W
R9tiEctcs/2Ql+mPevS2GT8GXY3iClzqu224QQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YO19p67aT24u6CNTYXEtxD0EjBQXNalxsdumuArZP9RZtZHyvN+Hnze5t/eeWwCTgmNJA555BFxL
Btud59tPSRiriPuNyug4aRzU5tot2yY6slFMmsv0xDYT3wkcNirJCgQfXRNBm3SCdbiGTgt5XYBB
lAzCrLkc/SWFYEv+Qnl70PP6qgzCSxxqMAQ3wh/pirdVNseL7msrTjYf1qB7so0f2taMf687uMbd
VF1XMLl/M2xLd4BUUJ0DVKHEhml6kMGd/jaDs9xIiWPBhfbtQ3znnOntMori1sokKNmycex84cTt
26NNAIikDLOx7hoe3D5yhR6s5WWSAB9QSKb2Zw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DyYbQFUgLMv4dZi0S0h7bRug9KLFz7ea2YtreZpG7RswJqhCdlfHsvhv17yDEYIun7JiBO8fl6C2
3vhQdC78NSSzlzFPO+ZntZ3HAmTqIwE8OMrfeMtybGtNaNGrSYRrP7DaN6venSxyinI4tYkUrcs9
c+u6s305LF4H2VwGZw+5vCUBjAa0r1YJrHJLCP4q/jY8Thfnsi4DOWDvQD/2h/AO+nYMWXSmc06s
dNdILPxUh1vTkIUXz+BHzObXaaaHLbRJ/vtbigIr3NDlAHUs4JpUO4hh67T5HmFxI/f3VZ3Os2Gs
vKjVQK+ZHGNRu8qZdJecFJ03Imih6s4TVtgSOw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OJm0IreRHOTo2lFi2O3wcRrr03NrF76wg2aNFZ7Zlgg3uww1nDb0nimbuLlRQ8jkqOiVU2NNsVEU
eNJOu1cfy8xx3ihppkygL6Y43JUug5SAY/nbZPXlDEh14u7ZoWQGQCZoUbcmdZSphNF2TixLvBIo
PPJ7+/tMVlnyxz4/ZCw=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VrOQuL2LwKAyF5p0DSKiGhoaQZDUpIBCXQMRzAhBcycFRtZ+56foGmX1NFlG5Gl6kfis8Tfnc4oG
v24kwBlMn8Q19tRAVhBcIsx5s/AkBJhUIzQFKtVEMvro1tVpF7kfGpk117wA3oms+BLMl8yn6fje
Q6BDWwzNPkE2w+cfLR6qxJIZe2bptTJVFtCanvtsMqb8NE9smt/pcEKe0McfzmYidPmqEKjsg1/K
X6LYvLfc9wN0zegA9PWiBNwO+YoAJzzjSRj3Q6Fy/CK4AYuLzD24RHdmZHSGJHChAS0bs9T9MjTZ
0L4fvRQFmPSsZUGnxxQbHsxqPOmY5WO9zrGk8g==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 610096)
`protect data_block
FE8F1hVw5eiP8KisWjGTrpNMohaEUdbRqHGeXg5Bn/1RC58dgV5ajMpXd0zyQ6Qk4OzaKcr1CfTt
4U3cRMUp61ql+bjf1KH65KAeFDPuwG/UMM5etHriaSEYrfzYMe4fmLxJQwODdnJJOLzxPRwwMADt
8axPlY6mOh+wvzqD/Ek4rpcBVZlFKKXcKyF6hLVMTum0EzPEkcivkYrfv7W4lPtU7+YnCXLdo56e
I+QWr6lWsDYTUs4I+J75AXQuF1ag6Pt3tzs48BPk+h4awqPU8vngMNb+8TB40ks4233MarTUntE2
vUPV5kOpEPQ9/07lyKxmJPvwHZ4UYABs4rsLpAyXu5uhlbiqRAaDdprMNnzMxY3kCt+eFUq5AJyc
UZzSWNRn1AZqqzh3xh8jApuHrAeITkp5K6clrjgVoCb2w6MxCeHzNOryia7Js+XOp+AH+9KqcJ49
yc5Cp+O7FdxgELjQAcjQWwrR9vHWGm+ysEdXH+rK1DzW11Fgu+/KliYWoKPWbO0RdfhTA5oaB/0v
jKRFsTpluPh0Z8WJ84TSYi7jhjc0rDZpTL9kiU5WGk0ZhPKwramOYYFAZkgAH6g5/IjUoJF3A7HX
RKsel6H94iblTxSy6stmeA+XkNbgBnph0zh4uGMd3BJDGhJa00Ou90D6oipcOdoQP7jzniuZrcWI
VVvYwUTlGRPCq4t9ORs8RUniEJUgQrYCrPamXcfE7I+3o0r9bDCpIc+ej9RfDTFcE5krQzYXQ6p7
2zVnkZtwIMf7/uxW7JcNI+rdPXOY5rPjirnMthpPnqogHpAZTGtrofwNw4JeXqD6nv+gAHxWF5Z0
KfaIPCQ7hye781k5v/lYtSbvunorJbRksVCOuWsMVAtnQxEk9PWv5qxrTio4srahyG8Q7wlG4B5N
l5UrcDhd9bYNn189SOX/5SFJ+gfdVrVe4E52PH9JsbQxtqfzbDDqSVbSM1oJOaS+INFG6Xeh5RfM
erMdHI/J0SgCF5rGkeeZtEpLvV+peOQ0seQvKPs6+Itfn5qhheJnDxR3KEuOD8al7x49CJiBBeek
B+41kajBA6WqRSgbYqapbGY5eIVutV5jQVSPFpdUPORtTYdqBpwKctbE2JA+XEHpcmap/FBPYcND
f3JHbbjg1NiXybi8hVtrs5iI7XKNcCNPNbZ6Vyt96e4GID1O97Bn8wTQ9X8alZewWhCyurfQCmw5
8ly0AIBISW/51t07K1Sc4sM2y6aQ76PH6p/J64Tq4DFjvTykkWiiieHFEuuAfCHMFkXejleHV+XE
+uo23E5wsfa6576pZgrvlj5MoChRH6ZL7u3SMSFh/vwi2L8sToYErAjaVY+X71waKsK2bMEIX5Lo
MUD08/61REHEXcIXzqko3wDG3Q/o1q0ym2CUsFlr1Cs66qDSPLegMNCm3Nc5ohSE6ykhBdZHcZ71
xMcqq5TGa9VNVzt1J55sE6tEfLlFTQ0agWyzNAQkaFcEtsfytwaUayWNpKko1E2Dh3TqiNSqBiIW
hkkZYcmwdA79kfHr4WFMJRK3sz7Oq75RSi8lairbasjRJMXkvr7r7tsKFEXcb7/Eojw9Bc7in2Pf
knVxUUp1iEyHdhCXD2VC1bKAMRGWBKCojAJKFuIeAVSWTaLWFwMrVDe0gU4OS2+UUUY3QWlNOnLz
gmGntAipxrmyVAdCJAWcNbxmz9eQF4g0VZQX+AppgxRFoptOW/OVJW99D9HntDljVzjffqf8wAu3
zTeYVc5pYv4CI1Hkp2FTbLpblqgeuB2lrkU00noEzATUclW1bjF8mJHhttDt8dMPo2HWaf9qKq/2
4hYjDZ+0iD/kWHegeG8fFxrNDP68/+4A0cCqJxgFp/YntrK4AebrtdnPUg87iZkzibhRn0r5hqcJ
hnxvTsiOmFU7Sdr7dbtwVANrDgzeE+XuY3fj0gDTlktCmyeCxuqQ/A7z/vhqhsybK8ypbvvDefHl
MzA9VwMxMRWeqqvtgo3+MHI7e+NAIwQD7QFZrG3p1dUlDImwKmv0GkjMKDiLJQ1h6blvHi7LNsPK
FvCb0hPt03lfIEiG3ALjLCAOnjLiIaUF0daMfpFCK8eD5b9v1pS5SReyPTKeY1LsGMVlHRdE93OU
j/XWTyTINQr0C1vhoTFuVaTeNjwZag+B1wzDOyXP1tfTRCyupUoe9j0EAITjsaQqyoFhkNONyrLv
CoXNxHj8P/u3NSBJOS2eGIOQb80JEIvC3/plreOiM9lg8d5ou0YRhTiRNE/M8+y9CFYeHzeRSre0
jXsN8wLxUafix9A0ekQe2ABtIsLxdp/vA7FaQvzWrtGre1NDBIs5HqAXwsCzH5VwWQQ7GW5BVtIG
1tOkDw5fnLwvk7AdfYrDbBuwaO9jnWy5DvyybtO1NoD08fgnrawT6RS0iKv5hohfbNePnuuwLd7V
WNKjw6rIhLnp+C8mqNQml5UqSXxAFu6MwrWUPzhlwwVHVG+yA0bDYYfnP077yVYZ5yO/eX+39ywq
y8ltZ73m7bW8jzdlrEBWUZT7MazjRzgvXzVwi6je/yqvst//7h1AhoCYClH0DjYIE4P9s12zdu+u
ipBOCgKnGnqsSY4FVRcFVMLsWci8XKL4izpyYL0pGmSQvuOunJz8NvWXKnOZ6A/6OnekRV/N+shK
EV7j00hzD9byQ0imaWUfUOW5DtMkDySvQrPsxmVsj31e47pL65rX9rQfPb4FquGCyq33o+OuwNAk
QjIWZSjNy4fCCkkeco9bS0EzhlfG/hGC/KHza029WjrXOxt6yk6WSCYSle0Vb9nh8gA5tvr/lfli
eg2RIW+73Q3ytErexSq7CNg8MMLmBA57O22E0zPG5BugyUQvsv5Ax6TKs8Ut6nxzbniUNFc5Wc+6
Gh1nOyTEwNYzIYebBel2r9ljPU1G1WG4wDby5hHkMyl/6gUeiRKPGqTOuUMcSpyZYUWYJIicv3RY
L17LM2IDL0DdyVvebHuNRDD7RaRlcuEo7zF+mAG/T9bsm1uMTAvXupT2UtYI2wpgYP+12H8hkn7O
bolQeK6AfATaca7A7iHvKU1vrp4nZBT8Nn3CerxQqbPmXpL4W11Y3He75LoztASpPfYVMzP5Yjd0
WVV/UaXNwW5drnNsblGm9U8g4aEILj7iggPAdGJ4pbGAKrKvVFTTJS44MmSofqErQl+2iN1mAxGe
bxnUqA0dK57X3EPMJnE36OtyalZ/kB+lRUwdm1SlbK2dnnRYQGqgIGEeJb6VExSdqy0nT7VJOH7e
b3M4DTSmRmOIxkzqlGcS/bvn1Ay05tQNB0bH+kuR+DBiw9G8infwE6vFRuS5Q2CxsdlN9RkhEvnm
utSiqTHw3UZiLpg8o6jNux0QhxHJdHjprdLGPSjB4lHpUSnFPoqcHwgJwbHkEmQznpl6DQaQwAJs
y22nynxYUuoQMr6vimBThUD1nQkdaY0jvTavo7SHqnn7tkt0ggJJfAdxy4TCDoQAaC9BOfhn6uxZ
wDeSz8Gjhhhi0nVzX4sQDv2YVpVuP982P7uI5wTZ9NKwASJEWdlDshd695cakxUhDQnRQ/iPURHi
gMEFbqUHCedsgsbOgi8B1PqhOZeKtI+u0vXNeCNJvZcXMoXG3tFKUHbxaxh+/p4HlvyNQ67O+9SD
LEZaeeMCKJqTgPPLRhdBJEKU2f+/n594e91OZaTpnDFBtF3/OxUpMKLAChV5NOUy4E/wO8RWqsmt
3EypsfXN2WRICxCW+qyO85PrSJGb4oqIN3PeVZvwX9OKfi+a0/AdVXvpCWoXzf1Y3J/iiiVWEPzB
Ixc1r0nL0xefLN3l2F2VqxBUWdi9vHaC1l9nB9dhgDvLG6K4GzKgNRrN3isngNIc2hXw2JMQn1zc
yvre0YYHxsnqJIo34J2YvfDKUmgqf7/dXedBmSBJ0xu7Qw9I0ZOTaid9PpcLub4JRUZg5cTXJpod
Dvm6uZiLCc8plVoAkhTu4lpWBGLpaosxwm0jHC9OlswKvNVQxyTuchOZA1OnQLGVgeIJo/MA9a13
3RD/7L+fKKYp7/9m5l9cUXQmLhyQTkyUZMlszoNMLsJT/W+tC1x6Dj8pveNViRRkiNc5wAlKU5gd
R2HvpUvFjL8n4RdGBwA4RfIc1YJAe/8b4+E7O+k9ScX/5+SzInyGCGjyWk9kkAVYRaReVKmbY/rQ
0ZTQ36Nz3XFk/qytleWJ31LmR9+nuZR4OeeOjcY/it3yVD/9bUUkKQbWmtwsJlHQPHoHXIgLb/vw
xu3ejDdNP1bpkllk3rXuNC0be6boKLRtsBOrYYKm4WvXNQjp/MW8eHHnPQO8aRigyONdOeLSlchp
DdbuPoH9L+QprooHFcleCiP979eLaNN9HWVJSWGBfq62n+b3tFEMQxFoQSxmdt4ylVpEtdfoTqcf
fqb1MMP2IysOawblj2B/eqHpCXbvPADMEB4/R2gxM2jPSlEZvIyIphLIAcXvqdyjzF+rTxj8BhMA
FWkynLGqeWILNFZ0UAAb+ea0Af/vjWglqb1+5uWtktHUEYUpN4xh3KsvGCXbFrHLtEgrFc6cflBk
Ee/Ozpp24kS4C+OkGeF+J0AcqJV3NoIqFBcVd71kRVPaeZgLB2y6znrrKTTyFYSp6Bw9tq5iW2rq
NvAScujaiOoUg3ufxMH4Njf2qV/mXuwJSZNdsfN1In/Z+ST0Qltj01U93SqfA5bOZcRqnkZgJDI1
a1F0GmluMv2dtfQuhdVhpDdteTCFpuV04lkiScsIBHoO/XZjwoKXN75dNSH+c8VUNHhyEVdwD9o+
LToXGNSiPkMaXRlAuPlVbw2TfK4A1XdsiwMVX6wcqdw6GNisFRLl00QhqNFx7stLiHWNM7dqfJF1
xCFAYlIOLsgwOtK6hld7ldmQbLTIloJyJ925I5QS7cbU5/oacowC0azgbTN4M3IgdQ2TVpEEz4Vb
Zai4RU126BEov5WV8esU5eudDtfLXuaMHg3LaAatw7upQEBB5lquQaROkgxaMBcm2kgOG6os5iMF
Yq7XCnYrqU9Zfb9QGPofCEl+9LzqgLuD9ao2icA1LJbIvQSU0onJgZrdGhD/C+6Fdh+9QgHIKGg2
+g/CeW07gSo2savb0Pw6OPaydQod4ErdNjTHgf+vNFW8ncJdmFjaK56zogsyx9iKc/M5vOj0mY7h
3UcLD/JE/ob/DUpUjpCHsbxJjuB5WHjW7wH0zH6tgWQJGObEtZSXFkZK+uGribJZjiscYDwyNiGt
aW9ytfeIW8YNukFPCg636oGxY+o1x31gX3zKOMbe6DpD3hs6BAZ/ThTDZeALVwqbnQ1fr1jrKsqH
nWBIiZiR16TU8fpwsoSySwvBFNGoGwZcDhB4QoSy9+FoQL5n1IZgvlve9SKKhFLn9pRVEriDPyf+
bKdSJ9DUnV6py73o79HtvNcX8zo1DTQ0mmXJsDa1tCjkx0L9rZxMi9Vlds+gOpvQ6v2ZUGjBvhk3
OfZbnkD+lsqVA0k3+zpAHFQNaoc42JJ6cqdOnjP+jRwu57wC/M0kRUW9UPS3eUf86wHEux6qkkGC
lKnvqaGoJO5Am7g6gme9TlQ6EkB0/Hyj+W5vpjjB894YRQnvWJkc7F/hezaUy6NxV4QAYZxx8i2o
sKsC4cQ07Z3ee1ZBpZ8h1ZzA0fwrHmiUxcDEZRH8esa8E+UI+TBK9dm8jkSxx5Zsj3OZ1bQ1rDv7
wTdbM9Yg3drt4aY7LLA28iKoGMU3UBtvbDHs3LMe9pAvLgXrcNWKODepvBvggXJg35RKba8JiJVY
d+xWHk7J2UQPQ4d4HSR75g6ZB+yfrJ2ssXzHCZ2Zre5AtxBDhnq/FWe2Sa09Kr/5bnVRx09qMCbI
zyzBR8z++PLtw+HsdsS731/dWB6IewptiH3zn18DER9fE8CxlwCGSYV0E635uXV5f0s9ft91X1Mf
6zYTdxy8GwxrtG1zEl6Td7w9h4qbRI9dFRObwpzueDsmeUIBlMI42OCzbnb2X7E3pnRs8eIVC+Ly
j4GuzC9MXQzBAPwyCDnR2F2o6k4N9olbW9IgA4so1pFKpDl3Bm0K/UApGxBIOLngU39p0VJJ0nio
/7YB0sQM6yHsnxYDO4aDA4Ph2pL6Jxio8/N/Q9UWKgRxVPR9by5Ka18pv/5j3XSN5AahFFyaKIo4
4+omRpUsMkGbSQm++KI/6w8aLgjE+Dy1ugZQesSLX3DLpHqu3L4maY4603/R8SpIkj70/3JJBjq9
9MU7WVn/lfbDgf+zMr3EiI6CNKE7Ytx1Gm7zGZNrFqatnsPlCJKxUpc+Ns/ygHCZOjlYfGEDVGza
ppA29/uClEU5X/+08OGlL/Q+fFWR0c8UX4NX5GEeFRxfvcbgqHueKopZNOPFpAaqH2sSmlpvMQmE
PuF6tuUs2lOC1A6kjcqj1E44YPm07qI4xbblZgwKPMCJP2FIR9c41cBN9wYA0NBrY35QW4Rb54i+
DJx6Kijmb7nAQDVYZeIZz/wx4qbfrOB5vp8dHfY9D8MDRn/KvdDNq6m1l7B6lWXCpgO5qc2Db8a+
FiJRdfZ2HXLaL3fqpWl4hpS1eXQbsA+d5CRkuwrd3igK9Ir5wpckatGwtmHysFKn1Zi/nNDeKXvb
Kja5JUIAVmBnkEwOHIk818Sw5IwtbvGSykxhOVHIeTMA2C/8Mk7Fc9NtUaBAviY+7WmjgVfvq3gF
irLaj1emqjvxocZMy1P1CYO2f2IALoXrAMpRMTcxBAEoRAaqzoKtzBy58l67ujRU/6BZTXt70GuZ
ncDV609YwMqKIFQ6xZhX7E2hfYi6I8Snd6FZk87xY+RZvtbAFehCebzitOtAPd2kGwbfV8J9DpaN
+gGyKVoQbX71s5K/mqwzDFzxd1bb+yULqdfkB7Aw9UAU9JzwEYvEq8ed8Pd9zNihot9eYoEdQIqq
WbgieH5C4tSyMJ605Uy6LzLHXU8WTBSXt/uQHNsO8gVQ6LT2Oq1WOtPVxBkywIiwrf1403DFCuS4
N4faHH6ACCF4sIIH9o7b5E8Rohg53ulSg2UL26hsgsYoYqrBN6DDuhbYVP/jfHHcQSiz6KCPr+9m
DxSYgMxn7wSMR3/OgAGMeLMiKKggnw1JpibRN8yTorZxGugTpQ6viXrXcC5pkXs+ljISw44OEF6n
X57MM1ep8RqcxgYAb/aTrSAbJR/GaNqCUuDHxLEHGcQLQ8GWUNhGbT0Y4a1YxK0NakamKXQCYCyA
5rXIX/jVeJdgGahysnps1lo4Lp/hjv6e4uliBUmqYhfEd+Qg8dLUQ7OxYp+lFsyXK/V67Xfq1hIW
BmLic/8r5CoyelBHH/QzgWFalIpz64XrGlTgB9bd3iPVEyHc90NoNIhe1hil+slPWc1GI+cZExnu
VUK9OChRBNypenB9cCHZyjTYGDT2/lUerKcQzCOP/sxIpkz3Z8luuolv1BhHv1G4GM8ABbIPQ4mz
sUfg8f5M2eMhm7yH+OHUZwR3PcNw0zx2PhRSnknGQLeP6VVsi0nGV1qQkjM0iLFSCvJ98rGR2Qkh
CIZRie3w1b/meY4dcvCQEbW8EDkqcc1OgexP3G8Lm454eWuO6x+FvjLNPpf9ub9MX0nAxFmqM/Rm
i4nbF0lQZ8ZfexK//1AhKKBEMKI0LnplRMfuFDx4V9P+ZomAPXi1mFOCfbcQDsyEmhuDugPcmWeI
ZTpFtnG8Xd/Cc7ZVXHUeOY7gWIGBlL1V+PjTkuV/ui0x6G0eJELFbNkFRwEvro+liS9/jZniE1bs
p9au7bSsrijicg/Uxhg0qvrIXyZ032LaLO7atolXGux6rIRIPUcKSQHLB9R+NrGglCGN5q1SlgA4
9fpvmk1JIc0Wy/AN8jNtV9mdh37WE7N9jdyo9e+AYCX4V/7xJtQU1RmbSqcrstqnXb+UiQ17n2+e
SFvUzx0vLCmxx31G7PwWlMVLriFcPIjzX55a3MqaU8/hR35NyciLfAIbc+Gig17RkJAAqH87xQl6
YIT3l9SBb6OfxvU4L6yZhFqiRWVC0tWJiWUCMWFTP3T6GL1cF2HXRp0dg4V66v9RemsZPRENiOMQ
BS4OMBmgX+fSSMXEXtx5AtUPEgaOdL/ZUO5AVI5HfoZcxRL3zlWztDPEA5i3QBKSZUkeRUMWRzg5
Yu0/4NGKsMGRnP0S5wo0bLjnxmwDW5KvPxHZuOjSyvE0CqUKuiV5XMuMQQz8TpdVPTtMbOqhTYtW
8Ndznkuyy0RlU2+QUgBP8PFBXypVTla+4u9My/3xkj/yvxFcpZxcb4wPO+D5W/q1/OoIseMKK5Jp
f6NCcb7i5+7RyC8Uak8USQOjfx9zJiyYj3+48f3LKSYx++S9VDiDLVFahQFAbaTaSvJ3RHN0uMIJ
OfMaFnzkWaJqZoY5kiFkcNZcE/I/hXJcArzTfhxmJKDafuPI8NOKBBR3T6kT5GIHYAzVOi4gT6m4
se8g9QBm62uv4LqJefDuFp7Wio1A4UuFKD36wJaJN+alz/OiivYl8b0Vc6dp9HWAs0wySZeuTfk5
ESfAut2Wp/5mA7yR8tjhosKkOF/dSllL2IknqoVZyt44+RqgESBjjjlIPdpbq/aOyuyKYh/FecT1
uwynDand4XdiROFIzovMAZu9UXNwW6UNX09wW/iz1JfwicpFLAamDl3LyKU9vcHoqJIBymIV1GPE
rqaLnnOePEQ+CT5Z9/15/9toOgWRPJc4LGshvO8WsYMeD5RDGy91A8L7zhFvlZcKRqQCnBm1i7vZ
kO7P01/l0XgQtexW+1/IayYIJPrhLLmZXXBWcnD5OzyUZcMQ6KfQnnwfa+hQSvNS4tbsrk7Gf8sf
we3EcTQzxeowb92gZz/LtJjqfPHlI+meejtRCw44/+9L9ZC722HxBNCYeyEDM4kLfUJ+HW8zbrwF
pQW9uB1z++dCreS+Lmoy/KAEiVg9sVAVh4LZm8Q5tPE/SIVlFej9KvmTM0/06r4R4PhC6L7OPhWq
g1d7TPM5ZoSrcXDVL8S8n9IHpbViTMbwpGL1fV4Ibf/A3hFBQ9Es26zEAZLgFlceukX9XffWPJTG
S+bZCDFins0RqqU1OeFWoFbJ0/rKBJjMl8ZtPoAt4jzZiykd5ZkglYv/CGM10TRs3Fmlkw6ywYX5
aLokAckzBaFwT5k5U3/MQ6e8PGrVu0X1xRqixVhHqQd1kfktsZDaXeogtXxA2iFtLjCN2VUTei6D
W7IpHEHO1zciz7veQyuDwUUQichV6k0KH8jB/e0rFDtJwOfp2suzNmGoTvHwUVc/nADXmQDmwWZb
/5dvk2qSG+iU3IVViuagupH8/vW96skQnTx+GvaOZtE4V86iRK2NFgOj7RBrLDJPEFTL5ooEZQtY
Nmey0aVtTLcQHvAD7/OAjZ7xgPaMEKlzZi6N5DoYQRoqlkMCHHJgUUO9lrUPN8PTTEls0SHeRQ1Z
spipQjHPsOkkcoQlTE7h4Pcz6mfT0uv3jrLHPi6vyWzGzpjbNHDe1yuEWjWE9JKg8UWPWy1RtKwc
gzEw83C0UhxeguTyYjTH1lOmn+TG1YJMNLBuTcHGQxsqLo2HOK436SXywCq/n3AUB23hfVywFG3P
hi5KW9bFaFSuKLGnTuJzXLk7X1fdh5IYpGpyZriE0VGm4UbdBaoCZ5lys1H3tNFPbXHrwx8HIFSQ
HrYYyVWQ0T5yQA7ePcBn5RG/F+1JP6Vjk7zgvRc7OWsFtIhSBT9SBCcHMkLfU92r7V0tqrdSKzeX
5Of6FjCsst5MfnVdzSk9CAmjc5TNdAFAen9Mx2xtE4eOl0dFcUKRYY0djGOsHOday6t0KpP2tXSM
JonE5QTgsW7v9CPlozY8s7P3UMRyecFBITCAjvHy3m4HthrUzgigUrQXlI2XGPZF41GmPony7+Yc
V8CEOt5RhWnGNfhm8P6yT3+RM2yj0n6CdC4Nz1G1pj6anCCnm14Kc0FkfpnyilTD2aFMi9lkpXV8
bfgC9VWRwhBjwQRXse/bZdL5zbrBlNYnYUPpvJ/OjPKqM6erUFynC5+tCw8DDKBnDIbUXJZaUPbc
MNbGyNpruH2QKDxOaPvtBoZG0YjhTkMZKW0O0ew6nUH0iiQvlz6JRmbsT0h/QOiZeZkyIHkG+opr
g6jVw0rAx21s+jEHHOn/mn87AILCwg6CffInNpAxbFKDNQhrtKoI3mVg3ADNcq/NHDjnFVK0FMAl
MkKuNJang254yqdDrQ8c7k4Hnxpj0mXE0l8fMRviqTY1P20dNDdb/W3ISlDJ6QVI850Y71MIdcdC
mAdI7Ri/fi0LOq2S7+qvKmOoaHWyUF/YKmuF3hHOso17Z+aZbEVXL4j4nrDMgov8cMmoHrPGiplU
W53DrgX8eqN1dWM6iwi5uxH74WHCJTxvAaoPdurIGx9Hw/8ZjYxRHMOfDtB70shgdv/UgQTGiGfO
xa+e0mwr0kkN30OtnbJzhZ2VQ26Jyf2JR9m01hxzpxTArkmqIinzf9MiNVAEbBuU0k9Y6pT51oRD
3ls23tjtYbY6PPV/LpJ7v9KKugipGkwCMIK8hsTRdSkPFXuEq+TcxQC7iNV9xYypY6bgKOh50Oku
tmY+M0I7tDT2MxbFYLVhdTBiWRQBLQafFiqnu7OZB5OHthESb9rETZSKBDq/xEg/IHmXuXnoI0cc
O3U3pwbsiR6jOPO6it9g/cC1w6ICw4WY5a7/uI1fP7rwwlH7zAmGUQu38YBk7F05Cqft6PfaY6RX
Mso7tX6ihiGHVLReOMDV/7w4gHEFTl65tATl+cFj7jga31cCmqbS7nY3tSKGZUvxcOzOKAftbhIQ
+rGwmVrEl0YDjdHICPxesP4jbWOckVSZ50nx9M86JwUly/KUCQfqbCSqh/4tTOi+mhxjM1nC5MmO
Nb9TipneZiKhdajZcMBMXE8sJQacR8p4+3BYbcbmx7lRCqE+aBuBipZwziUffdMaI4PIxZAfoX2T
wlC1PiV8e8RfLVBF5o7o492LIfNaCErxXwqK7fpxhOVO5sn7ASSMRa6pIVNduc09PErRHC7d5n3q
EeYcGIz9qRt6XZlTvrUjV4OjQLH2bDHCPpvL/lNrZoeqCk/233Px7FLSSXlQ3Y5tlnjId1c0pCuX
MZnC6IpGVjKWJGucBRj7We8uEc9ntmBP1KL5nVwEYvQrG9byPIgjx2a/pXdAODgFzm4rAsLzZbLM
0pcFlqhZWc90Ly8SWJ6oaFam6Jec3irE0BKYSy3NLyjODcCM7Yi921RkhY1RRXC3enbSojOhED12
LcGFCUdfCn/BJ1zVgWqNDM9F4vm6+NXlbZEmuT8VQjtSiWbGMzXt2IUbg2shEHjQhn3chK7WA0Gn
AuSnopXmYin341mx6Bl2lYD6OPIvQUe6K7uLC0Li4wRusaggYnhz02SrWGtLeEnsKmQqw98rC10P
4/eq+T79xrWDRP9GByHtEbQEPIwawQFhldpP6xus0iZTbwbNtyoBIeH9VUrm+TsGFyDH50LZLm6F
Pah5kd7ZaGQIBj2sbyTH9RfBWnFoU0Z+n5hpgN88A83Ge1B69hLMJZBDi9ORfbJl/HWN3R7X27bW
3lzpNTDYhxOtKUhPoP4I9V1i22g9XhXFBJpqHak75u0yyzmw1OUjLHORmkJl96T02hF2N0IBGPvJ
8KdukNTC7XsYo7a2jBer9Z0Wwbi1Mc2L+3lLG+oVHJ+oa+tEdG9epoixXOduFN7yBHd3m5zpFxSm
00rE6c8KwwNGqcfcc+9oFsN/rEP/vSdEHl33+LENIOb04Jt30q7OpK5hMNRurCXWPxEH0fD3LSUb
OArdSTzJ+cyD2bSx6/cPHV7r5NwLBQNmrfxdFe0BLryOmMKtbvq5NhVQvuXRHSps1lOc/vbVxZZl
P9fjndN+Gf6spMrKWkmEq2MEigoiKfFwO5GlihggHm+0EvX3FlUYU1Iwee0WL01Zw8XSOidEJ8iO
x8e2X+/QgDwHx6bHiQeJBSS+07zflxRr8qyqwRqJHRW78nta+uiEMBkJky++T7yuszn8Zai9LciO
h9x3xPKJ2jX0IZNfUkZ+u1YxL2IkWppqVvLQp6nxububLFpzTQxW+fJWsTJTxyfUR396dS0T6+Pj
aDhupojlDm2bIEFKZVq6oeM6/csdzuzx8Kr2CSmpkpm1mj08QENern0EbDh99MWTVVFPw254ou84
V6FV1N52xAOkFymllnk6tmOlUQLpSDNyZv/I8BvOXzWQAuBV2OFWPGaLC4IBTryQhotxvblqKl1b
XlbdS/GTe8CzU6YsnQp2ekjo5NMCscazQz3YEpZ5H82aAivYxRyqXvqOxYy86xeOxzMkXSZDszBM
JE+dFzfSAo7fPyYtYDrtKencZqiZ8h5FwbZOKVafEYwc/gJXMrvxRTjJzoqr99DTgAQDmIs4YohC
ukqLnJp56bl006kSmfeTO6Wveja+wLWLkJIJmAsyLspb1dq3TEpHmP0IpI2GSebdIE+lLe/RlA2F
KYKgmsevVMScr4p6B3tnQ+Z+G7JebvYAW4JuI8iYmnVVQK1Ui0cjhJk/sPlT/tvtKjbBOItMkGaj
JSy6gqouq3r7JrEu/BUzYPhGgzd6m7zVyMWlteLJokuSi43CB6cPHuIwaSUN21O2NQR0v8RR8fct
hxKzq1YknBcYeozVeuPN1W4FlOlmU3HN60RTYq5F/v+48jpkpR0UjRomhDzqV0QyAGzqHTAWstzd
4pegPyzhSwDTeFvEfuObTzXd7zY70jq+VBTnmox3on5iu8fqSE8w2UH28cUQyAA8cRX1yxFbfXdS
eyslNz/Jm/nudEA4jlHTDlN4mRIY6LxGTmFG4IRjVu0/jUMDdG/kcj4rXh5STlvoP6PNUIQL5LKc
fcqnbyDRnvZ2Jurm+vMa6+5MYFq18zFwv6l/5tZ5fHqdlCXDed2fBURRD2yoIRVNhj7kwXGPMwwI
Gy/XeHmk0aDMMQmYLDh7+F5eglUAnAoTjVsJEg47Jth5S6ist1OG0cjPmKXKi/sTTjBPhwgZNM+j
pVWpo2ujuQXLQ9gooQB5SMVz019BLcZSq7Cgyqzot+EzyVC4j0aHA/QQ4VQ2yMNiRRrH2/KEXpU/
GjfeNArFEBzM7a5B0SklcdXpE03yPbvjTfVJGOvZJt66gsMzBTE2YnmXNp4M/BjMlSX0SEnw88kH
kSgxfibOZ3vZRBmXWu7fXF8flDlV4EcK+832b8/6xqrWiTnLgIr+OJQIyiLzQg50Z+sD9r7vo2I4
LAqlP7hnGZy4+T1326j7dK8iA32h3CjgOWQZceLDYjn8dhlgEEPugXEAwIC7xzvzxrk6/MvXLmJK
UCLjjxsAo0JGcM9pC/x66J9x+1QMoJE1r63FN+fVXxPZORhC3EOyp+XsU+nXttnmIPk90U25Feye
WlETlqiajRaJoFn45st+mAILtN/zLUmymq5QUCQ0dkX8ZYvJP2XaGe79gct3akBdnq1JCzG4y9Jq
x404606tCzHOof6umaY6tAdDkuK3KFPwkyoNaG+lRvCnb1bZzulQwueqe+DAHd5hAeGR11l5Hw1e
ca/epClhl/9J0wKzSlHJZtWm8ODZsfDncWTgzCVaVrvj4BR18naOOXuJBtiEzp06C0CkPlZ5T57y
Kx3YjK8fcc5X3VbD9xImSZxyRSIMN8NaNDPLs7db4ILSc5U7VCshV8ly5puwl1x2zoGJbxgakXER
ShUXUZeS71UMkFw4tLt5nEMzwgGXWfdAo/EjFf7qyvpcN68WCgKN1ti1vIprUzJAjbgca0Gktu9c
OVFFGfcLqFibm5cyR2MmQCc4mXKJhqB3mlFrkK+bF8U7yEr+BU4nyRNx8uRdMjpgdu8CeO2fSdNB
wzsInMrhG3b7xIrPkjVN8mNTq2q02VZtIhhByTOOff0rQO1JjuhcedY02rVREegcWLxKgAL8edh2
zdfsriVpl4M4uy1HmFbRubTIuAID0yAzQGphVDt7hpfOMB/A6xXJT2MOIYvSi9Ue6lX1VAy97++g
dTFZPkRGqexqHNb/jTbBXdXqWaJNze2diB7f0HZkTKQVXLqYlvA+lSPnFj6r5isitbUHbUANUdYT
v6RLp4BcQCtsUyI+C7arj/5yx3zUVHOMs8iXg1XVC8M/Rp8GwB3be3S4wlayCGcEKwZHrpsI7Gbt
tsi1JpkUCrieltwG9JOUNbrDpnu/vGdq8LhlyagS1Kx+jOragJP/90PzK8jglhiV8uRB8My6ZkcQ
Dtw2gDREwQpVMU5KhrKUF5leWKdPkJWfZgMDNvMcBklpNzdNVQwEVtSZ8ZL7yWU32igMrpQffkaE
bdSIlvIz7ZFWlS4I5XRHpI94ZarNpyhVIVpsr9fzCPeozCYHxlZI8N5qyzkrh6OZod4979KOEhiD
4PEXe+bo5vjOzFmHHWji8DH+4coshYLT8Hqw8NfbCoEswzSC/3Ua2960oow1X+M2vP0UzGJHsmbD
fZTsdxxlvuFBrHRcWwD7FhfUFd6Us72asM0NFxIZ+bXBsFgw0upPNuKJVkA2FaLkt9BaXJeany16
ScodqgZffeViUipp0FZmPrrpv5q1smQb6Smzkrum27DTr70bXS7h5vAolbMWHVUFPWN72tSBA2IF
gihmWg0PYkls67IhHCdL4FcGWs5QYe9hxYp6AUH0b/cO+4Cr6QcDiSrlIbF4clIHz1D4c+3aBOX8
IdGVimex6EUqFonbC82BO9H6g8Omr6vu0/sIaSXOQi7dOZbuxw99a++llnnRXH17gtAI4K/Ex4HC
SraHQLFqykNf5hXmWJHI5n18/Ld3nLF62jV78rH9pEkcppR8mhXNsrEAcldq+vlHCwNilGlVhJdW
BSaQe/8hWjs49HLVGXJKt8bmgzvI6nDjfpZRtmTyqg7oTChJgto3tY4N5Pyyq4Qe5jZ9qVBwJjw5
h/z+3mUDU7RmpEq89iv9QGCKeReRCoB6Nz8mEcEn4P078hRvLcP1whBOq3eSdrMP60IUDobng7RV
ByTXWJNaZkRlRoZtZcQMQpeisBCXdbyjtNvDOrXhYnWc0CZycJuc6FNRA8NMLOLUzqIq3PsK1AIX
7BYEcCQ4+nANv0wduQZGh9QrlDWlkUkfiEnZHKjS5ERFqVpSVxOC14dz8FW4aLLJ2HJiu41Mj/jO
5FVZaniTo/G36c/RXeFUEEQ/nJLuP16ZN+9JOC1LTS3OHhsIp7a2XYHuFWl1qCchK9Txfu7urWeu
bNMEO/Jmlp4460LJk08QAU3sI+XFQ4yYa0xXQW/PQHbf31YuQ6WyqzQ5aS0G9/9gFS2zXaUaIpuW
FxUobDopA2LBJnfX5AEdOIxjRL6yAVhN6UAkw0jhbafomPlg7VNMUmTy7rjK3OMovcUhow8dcZJq
0d1TgdEp+JIw6UiGGFdA4LZI8CZ/yTFbpZo6PlZrJ7a8upRW5qFZ7lv6f6hezv0L1e5n50cpT2In
VKZFBeAagDmUf1aphxvcg88DkoFA0Icrrumyr1yrUPVRbYeUoEuzD3bw96lL75p/DnvuRQcxnfvP
sbM6Hbh371sMpeP5+cCi+GPUXHxmuw8FzJQnto5YSlIAF08LC3RHGlGydoiheSGT8HOJUSeDvwtj
D0tZaB4s6CKyoZngVenwGs1zb5YmW6oCWIjZsbPNUJHxVhzVB+AJaY1te7aHjcm0qstfNYN0I2u3
EYVTedG6W29mRTI9hH2zURV/Vm6rApsV12oIOQaKMqMiA4VvO0KqeNHJTsQl76x+fD39q/xG+Uo3
IvmhfwEczRIAlm4FhqCKCw5DY/LKJFCN3AtAM4GvFaClb92qCdcnInRD2u1CfCKDagXUbj2MFRI3
r3jWvPL8rC1rECNuyBXjurEXyDEf8UnyABoAIbxw3YVTIQFnjPBQcNnL7WjynByNK9HJZuCjqjVr
rXJu1nEIlWx0oWCr6d8LA88PJx2D6IjC28nVR5L1iC4abWwYX5gfy0prHfOeg/Xhcy7J4f+pYyvV
ctBpFtCyob/5jnmDznFXIUG/az/4ANHQFuA0zVBiSz1x6Bl7Okga2AKbk9Y5jzHBfQ6IRtbdxqBB
nEtd7yqNn0kGeH3oEmcP9rBbTHyuky0ZZhqU23dnFqZy9UWlvdjQC4V0e9cChd/+jQLY1yDi88pJ
93OwYiGTwmdnMAjyt8WvViLCZ01nQNM2bFeYE4i9RJOUQKlaXZfQ7BGFDib/DXFSKNrjALLnACAx
jw4f+xH6vpsFQrMnNqX67qi0m3mEuwtouQZa6wHZRsgEy1AMk8XQxs+bbo3x4PBLXHf7SC7omoX+
DzJUCcJ5uqeFxnT4w9QhGNQM+irY+QgXHdc6fk8Wy3CTmpPkB7JqNdp4d6r0HSASe+qs/ujd7oaH
r9ItBerxY0K8fPS/pGnZc80XC3cRPW3kabLkDsGRBRg5cx1b5wQ3ZldyXZCkAvTV/Dnp/fAbZhvh
73Kvgp46RHMgx3/D/JQPpPZgJpSGfLgFS+FZmExPT+4AQ2Ety0zv88VpbmAwYRTf+OVAcwYgM67F
7N2n8WD3H20pyyVU26EEoI6s3AhUkF9Y08u9c+4JzZ4vyqdj3Hr/yKLqxT77faEkl4cl/+A6ediy
P38FfONuHsB4vZ7hWPsc0D/TkIQSrXjfuhKABe9LQPmHbnfRGNMAJAS6YCxei5xcjJY1h0Fzl09G
ocD/oV4njWYzJH5khWrI6VdYrYIh9ctu9owXXzq2xj7z8vewOy/tmuvMax9H71xTBQ2N8rcI3s/P
PgTtFY1T7fkbaNdUt3xIX7OWJ66jOYi05wPxXYiiJYuY/SMiUW6GEwE9jHG5MaJ6usFascY8ug/D
pgEVp8Yu6ErnlPoy8vWyoA+OqRqKWUKQCYTOEmuMuV5XhaFtrnDCI+FQ5BFjHg8WHGX7uBeoaKD8
aSdtGsR+MR7VD9SiwANxe/dgPZto+4MSJXqSIM8w6JTyS9WT06WeK8PZiTWAVzq4IL44vdvhBVrY
zNJAguDuJIZr0gv7BWjVS3TNuf/6wNPA7GCotVWSOt1B72U0DVW+o2Q+HNdWXqY1VlJ9NGJABhe5
D8e8KCGU3S7OYell0fvqRW2UsYO0egit3iWzDAyg/ZjeNbcZ6fgTIioXvexHsvpwAo0MhGbN+8MB
mEIsAT5NOQa0CVrSdZXGOBYhAyTEXIdW1JYjGHy6eBIO+XnDYwLV3ADgomk9pVa+l/JlaiAqdNiI
JNMSLjJy6rST8dMOWgzSba0NxQUICzaQ3Y7ERxofKnMAXdp2KHGaGQVyI5kT2IZCdUBZdjV6Iily
LWWISiUMNHK+ThdVWldsliKFQHDFah1ZLQciWQeqG774eayXlEN3syg8RmeWhSEKq9QpnVtjr458
mXWUZ/qS8t1hLDeIvCQZwlnmOrORoq8yJHBO3CxSfy+Ih68IT/co6bs9AgqlGIEmANy3/xn75QI+
tiNNMw84+upmINDBqB/7ZFuP8IAmD4/OfIluJRiYEBcM4hYZ/BIjg24j7toyyxf1Ai6Xz3qOpred
tVTb16ZWmBDmqdBbs45WhONbMzdQdXirceFNKKpZN191fAKsxi3y0JNXvihiy8fibVoVM8HR3ePq
BN2GBHXzLzYBMihR7ro2siu+snWmLn2YLg/ZW6X1Wu3pZoPggY1d3PCPMVVmL7K80rJuEQqtP6yB
so6wAwo/oz72JLZIvSEA79sg4DMCKSN0g9OlQsKKGJZkYXySBXdTPAmMQyYoOG7aDw2PfVpMazSt
Qi4kop9nAYlAcf3R77R4/KfHTyCUm+ZELds9woYWzleQoTpmnRnRUBqND7mg5KAtRgJe4mVxgR+V
W12DQEc4GY3FBWKiYHBbwkZcyezpsk4YkXz4zC88sEC1lqAK7Cs0hETHge4kUc5TP0kS3QGr0j74
vXcByEG+8wkbYuommSqyp/t64ptakDt8Zz+jh0Mxuip2dL24GjHb1yPMHzkQC+UFskxmqA14Qk91
5b0+m19vkfWYXehqB/pKel3KyJMoHFybPYXE5WOpdEPnLlRt38e53Xzg3EeO3O6JKD1DD4QTZDPn
SQXFPzzsl+ZwidObaFOXcWL6KtGk1LyPQcAn/RAOts4HfVYh37oHP8wVG3IZMAwYjYwo3LWBJ9DZ
alP+BptMqZCwuLAohd8K6aSu/18H2E3QWr+2xptQkFr9KpnWtXlcY9VNW23Jiwlawp3NWj1OtoyU
sl8Y42ypwsFramJG+kqiRtkQUeOEqOgHzJPORPc4/zVyv3rzP2u3NHx/VnVmDI6BJePotfxtb+nV
Pj8TXJA6vRajCiD5KfmavFFFBRoL0QHzCLokFN82Ap9hgfsZpJtY+i9P/h225mMnqNhbD3rF2gfr
uDcgk9gxi6ChPDH+XlbshDhvbKLBKrFuv97qP0dmNjfGGbvxCxA/u4pXLgwghPhYl5kOEZDTL0SN
unfBl3RjK9GTznrlNjk0RiOExA8DvTxMZQcyYA9OdtP9WhnM3p4I1WYR3Uj44HdJKZSuaVOdA6QR
o0CcOv5cSgUM2iyiA7SOVyKfHzD0sUszqSbENhO8exJKuxiLM5OXCDKVA7pVH/3shnaxLOmHmd/g
M+8zEGnvs4JXRUyE5vkSjvWyaPp/uJ6PqY8+KRAmp6egCDaS6c+clwxHk/vRSG0Ts6bjfUOXOKxp
9YLav9XZCBSjkqE4OtEr/HWTOkZxC61ebXdX3YtZWqY723k13p1ElpIe5oXxGQ6kUiIfzMjFnMTl
hodlSpiYXhFgAKxsZbC0VfzcnSQ5Milafzr396OCBrlEuQHqk4wLhbmIqVigUkFfV5ClqItY2t/A
qGrbvR6A1BxEiu+yF4bB4FKebYNyb9JkzQm/fCQeKtsxcR25pPpX6WM5mOXbIZd+YW8fwehc14fW
kz8rRw3JtqyXVE9kFSNJBfG60OEHxf02EdIph7Z0mU+lpxyvSGu5bBfsyc+CszoBQYHI2VS2+i5i
eqsWSTvXR1aNkjFCl5n6RQr8A9ac8MoXhDz1wYtDYk/H5qJQe+FRWKzF64nOKf8wxkJYwPGd8LFf
g0LMHlNfXqID6n8FAEtRBejzWMegsEMum8BfXlMwuwKOs7GXpUPis/yO8Y/ckIEPYOiBjOwdrqfY
51vjmP+0JDC7LeTz7H3dZhq+NR/n2155flwtHP6eaVQ6UIZ8H28zDjOmjrIkEHN90XQ8q6f7+YjL
VaT4ZZS6TBX3FnNGgBN3O4ZGjn/QBbxM2zMbENOX7FIstPxZNrWUTG3VoZ/rZ/Jmr8ov8LJPcrKM
ioO3i0+Y/w9+bPAHJ4mQawWECa5mYRekwlywfEFjmSVLhRo5TO4SSffwLTsVSUO09Pfrk9VMGmP0
PtU9s0hrMqM64pEKIFXbmPy/0xT9IFb1Xr8NB3hOOcNLUzIpwbeyuTN/IeOXim3rO92bK/MQR9/2
f6giGiLz0Jqcb8QV7h69CPWWQJPNxdLljf0o/XJgGhoei1aUI7h/1AxT7P9dBNIDY43PF6BUxePy
64BwYeOHtTqtGSxQKAoZ0mzSqCZjNa8c6cfDm1WGAqkbNLH3X0xj6m58frfaKMt+6XwzR3LblC3y
W0ipl3XylXABKwlQK41Ok0qayGoQnCU1ZvdMPjiZ+L09KMdP4ptQJfofCaTUJKpkye2z3CokPoHu
kdrsGrcOkSZq1yrJM7arfJUFhVSnm21EEqX2jF/D14W1DU2yRUNcDxjfRHNVLHbZ3jYpUfEJMqD8
3bYh/KRHsLP4fPPWG8sdLfDEqHKd9SuNtFPMD4uwA4kLvmdAS/w0ymjXrw61eXyK5xaMR+VMrnu1
rD6snzD7UdIxRvUBUFxiRMEipMQSnKsN1YSwdqGB9AXvz2OefK9JL2mJCfVYlwxb+bUnFc//z0bN
lPaS8Lbkxm4loKmvqY7bj9GYci8mTvl9MiNsfgG/P1/grnrU9np41Cfa43CvznjClIP1fobLxrIF
Dj3xTC11RSQpnUQ2P5z4MriupnL/dDNZsjTL47fdjHvHadQszgztiW6IijoeMnhTnq8tOZaNIM3G
jFWxg/uJg3qoaPGBsbucjZofeC9HkKpMZY9fWrDv7G8aHt+UE6mihx1Pb8WokXanibVLHtvVOgL0
QvWxJDJ3JGFv/QuxqCditSeSbMPrNiEcx//5nK3f3E+qS95fSKDcwVEcVXW3i7oAyS9tvAb/8DFq
zLLcujuvDyqbR4nj+4CUy+zQEESJpOw5BkEvdNjgNNZqyYVK6JmcZ47r4wly0KXylzzshnuRlbrF
Su9szzIHs/ZLm69gNVw5po0DyfJrO6ki6zCzTupNA8wMdpezmQDi78UR/e0ERMUFJWoAM7ykC/cY
AK+hbMaX8x5j8JBZp9tsX/Rzb8ZwGUE323kghNHfq9SzqEbjQz6/q329M9a50Tz8CO46NIFfK0VA
gvRfoLoU6LvPwFlUbKnFLbkg89jerbkpKY5nMde1jNYam++CDFW00kW37DaxUO5hldSZJiBghDps
gcTlim6CRkZpNhlr0F9T3eiSbsWA0lyGmMpfjsonAkXzPq8+abQTCmJuT8vdNGxI8V4SuoUUitPg
VVPRnEllbZz9aLch4OYPFy8+qUBPdwchbNaKWddolIm5fQxxsswhq8mw7wGPGRsnJnnUNXjL9Vuf
FCrkqV3tRgs4urk0RpkMJuujorW3G09KENMhZLMIk5yD7JxoYNxfYjzJ/NSJRpgDZcgSGUkGy6ed
ngCGu52RwLPRxZt+87IF1cQOCUrqUdMB/Kn2pUSOEJAKKnxxZkBJzUzlgTlyDGBTkPmVORKOEDnT
0VJzgcryeb8uRitl5KUcAlpjRbN3++LdhAPXdJHV7drxduNwfsx7+T9/Li6LDmij5xjmQTWyDw99
C7TmjQT/3kU7myHAiZRyYzY47eXXYEy2KX7LjDC5f1Owpl+yw2EbYqiTK/nIlCUPDsGLgguVi1SR
L3JeBevkc8DyzREx5UL4E0vVpV/qifvFwEIYdcX5ZjXBqylZhfAiR8z4DZ/48XHDIJueGmrlxN0V
9XTGlt9c/hlr3oK2qru3TtkvxgdJDKLGmS8C9x+PEp9V1jOq9CjRvUtQUkG8E4hhngpcWJmwdJkf
iBR2U6pgg1Oe4w3ctO1XMO0yD4CBCoYO1heEom32X0ZZcfb173oOTgIAkNJ4siveSqF+kQ9GY5Ni
kaAI04HAD7tk/AoiHo5yc7bEVaRpThEROoTuwl47Aec+BKBkd8/7Pes9GoL9qyEoDzrUp3NIfLbx
bxQlfO+xyM5k5W4DaIW6KvkkRYgyvosshYwEvOQkLPJNx1sQrS9HVzM0/8s+heiJb+pCLRzs/6dk
zYd5AdIcGKCgnRszcqjoT4S9kNdVz8cpy1zXwdVTnMRaXUa05/ApZF909vgMrRbCtPUJHaroLu5w
r79Di+dMhFbS8/qrSRLTVYG4p4xMRNfkewGOQpqeFeZEZgb0NYBsKtDM+DNZL1GfV84il1dENs+J
+Ahnz8VPHdX6ONQS2X6Ve1+m3f0YYi3RGcohvixJi6DnQC+WqmvafkpCuEGtp0NCZ9AtvwE0rryl
TANcLi/tu5B4qlxaljJ4cqPSdTb3EzG60SRm4RX0JhbAK50hKvUY3aT9atz9zqBm5gcXOVNB/AQJ
4rsNqgsDkti/E/3SjoDT/x0gpvdho87a6zqjjIf8ywhPlrLSLr0DrPa9XlRDJD8cxLonbxjNRYKf
EFJrr9zyNiPj8/3M/5s3WH0q7PmAUCE/LZ/Q5v/9RqoHhGBqXdMG46ABQgodVwicQicpd8HlULQs
LAEDmNiF6yYkNipLgAmY9GMDU5+CwA0gbrPvHuNBRlC4ADmiEGz2yYuvs+uz79Ss/CHxjUu9oyFo
GTEEESi9bD+WmFBUmDstN6ad50bAZd034cgEJ5d88MLinLeOv7hZijAxMYCGFS+Jk9hzGlF8vY4w
wEuHz0a4bHG9YVHMzAiY6lXw/lXMMd2dXvCm56QydqsShD4xsxFUr5on/2p3YL7K7uNse4iXINgP
Lw8UAqxo14D8ye/hMVBTd3ra4mOUYiHORIO/sg7/iwvV4sP1l45GEqdxIR8+RdIPHR/iQomIkLg3
NdjsLhqqTcWW3LbrqJ7KzxPFq/+Hi+EP1mWbbG+tB+TydD2MfAZ/WLIyOxfhoCMRKhefxY3Nscvl
imWq76mWFIc4xSXAMMJMxpyOcdICRWXAMT+FFpYZA5Z/+YOoo205EBmGXRm5RJ9wGZQR9619lJbE
BJvnaJ4+WEem5ULDVC+8um73MJ7p+0fF/owdzDofwPX5baMvPz8P9lbht1lfbpXY3QCZNLuwDzdy
YJt1g7LBmHOX/BjB+0wFIt6fgAA/HKH+6T1oln+sMIkmPMZTGEcYoWSAICKyk8wJ9pQCjaJEstgy
d5Vc4/5Hc9+sL9R+s/E/W7pB/ccgim12jXN+OJCOi7vf6Fv+zA5BhpbFQxjUEVIQyh7XOtd8bqVi
3Z4xVhsMP1/JaCGLLE5oxgdLTMS5M8QdAI/HOI2fJsozqrWNyp8LQAKE63+3K2/tcXt7x2cQdvHi
Nb1BBk5xEAtk/FS+wIjD+m/1k2rK3XfsgiXikLmQSitUb5PNDXX7i+FkzXtdcrGEjdx/B2t+UNSN
FA+dIo5iM0NtPFrIVaEaXjPaeVlWN7lZTDJxKeJlnTHddpYDVQ0m8VHNF85hXFbZJnknOwn+m470
cSuerbb5L6fKopJxTA3htWJSRu0Plk45BxmWeD1IQHVYq5Q0Qa3cggZ7VO1dk2+ukGVRIEW/8Ll7
3+n28Yc4RxlGItTAPy1a09tnh38ZGveESCHn1FfUSTcuUgsZ9Y7F9v46nmQOOpcEXIRVkk5vCNfQ
RKMLvdlt3ett4k4LTPyUBx6z5uMZ2VwhA9MsRBgV7HpZhfQ8vTe5ly/qeuSKgQCBQaiiKHcNQJnd
VcVtoTGjr+83WqYFlodYvba7OSMNu4k9OWCtR2hCb76lcv1KRbqZwR5DlRe8ahekzKg2vdR9RH4V
ii8fdxZUpkPin7JTSuyplnyu/6KdF7u7VNO0KR5n21vopXv2eLcWRUlzeAXYX2BrlpTuc1Ifehti
FFQnzfh0UycvqpgsgyQ/dfN8fWfngid9qPoVkPS5NZsZQJRhoRPHcPiSfxLV0jUeVBZk+zMSDcC1
lJ+Vtk43ymMZTPqO+YEC2wK+ao9lZN7dncOWofWpPNjEqnkFT2sHupcwTIu6lbJiTqxYsRcQvEgq
ZSPunMGw5juWLCplTca3zMPLAoKwRpal1GEnfbPtXHGiStt4BmiIdZJ2164JI24cfu/Sf+RNFhH4
lWGm9ZZ52TKbOdtm3c80JKY8wpdSK2vylBlVIsLs5aonRvV3DwVEC+YsJCLHuSEt7RiWqZb0NqhL
WP4FlKMYqyhtIMAsIT46Eeof2ppl3evYmCCmm2GfQNEK1UnHnRn1ZpaTBedW1bcVTYCn7x3YDgt2
788gCkmFmXlgeF7oITiQneecmQtaXYAPk79cT7y7zl+x+mGz04LNZFUDslnNOec0Z7q/z2+6MEjY
nDRoqY+PCEXnKaYa3gaDCFvQU4Lp9T0prwmuWoas382IwnSQY0PYz/oZLsXQ7MjuCXHK2NC01lhV
C6MSqlOXWqRYLd/GkUwwSbiVMDE63fHI5oge9WJqAhtoYEwqcW32nnabKsKngcxwMxBz4gOl5o87
UJXi/mVY+olNLcG6Do/UMczwDFcjSihEWA1MIebI7YYgak7CUw1K6pb94YtWK6i+4Pn+YQj18r6/
GwqWXCXmFKNPZfjMYYPJMMZwOrHK/O6Lweib5jGR2q//Jbu4fJdeSfwNICUcD/1QaeI8kumO3vWT
MZcCLdgROX6ZwscX34wCbVsY85RK7h1XopRyTUej1aeBRFE9Av2oODJX/4TqLSQA1azNZnpAKZjT
OYQjafx9UIOzeLOUHGqMi/r3TVyYpiTUEx2YLuYGxRzSxjBxWZpo08Y0oxZPtLfuxrxxe4TNuTxJ
dmSp+u5mfL2yQqvW1gn+VQxRvjHGejOWl3BPM6GzLIZR81RGM7EmC2q11LWHPNPYDmFzG3j+QKOT
idbn/oJBaZxG2Q7Y7JP5N4nIc2aLQvt8fMd+87d4ZcS8P60ezQzTK2fKBxQVKtNJIVy3ZpG1mpDV
3AyplNi6EOqrsKTbsG7+Bw+HqoaiDZOvD700PNitoREOYsyylk8o9vEgN3bBWHYQGcWZ6IGOFsRV
ylsPBKsghh0Qr6lvIxXqpA5FJAZ5jTymqXTdFsemko2ikBjulN00JfVFUbCYuqn09ssxs+PnqwUM
26NJFjjIOBEvhBxW93uXXkdkaEpXmsCIBwrr3bvQhYpA381F0w6JXLTSkmhYY3jUVGQtC+Rclz7d
/AZrAabe5De02x+4wSzu7cOMDbW9R4nbWMPizfm8WQiCtOD6pXTSCnjDLSPo6N63kGv5cIvSCj73
oUyQzgHlxTI/IL9vgBYTZVGjpE1KISBVfXM/vxCdFvzvbnMv22iJmNedDrbCkt8fhNb2yve4/U6X
DemwGiDt2AwFdTrL2fe81CCgH0KendsSFMktwJIcoBm3sBv0P/mvcPZ3fp0XjZfHMzr3bb2zGzt3
DZfg4JvflNWpUKUH6ADyKLHQy7wl+PxNgElYoVovjp9LhgM9LpIKATorT2sam0NfuUP3+yaCF+c9
IJNoPSoO0xjztyr0Z6ncqNkKa6Je5vKHkFvlP17C9fHW8WmIL4JKnewds9yQ2xUCL9WPpV9Iy8+S
8QHDbgz/zgjeMlEdS3udXdZqm0lhtupPfHO4SFfyt6K2S+t5t2Ony/zq9N6DFRJjwuOzkppZSTK3
MbQP+npR/UQukWACB8QSfUzPF4FKwaZxYA5PuGhFN/eYYnYa+ZRnFS7tU9MXGZUjH59wr/F6iLmh
zz769Qv+wV5CIe5Y1C3I4uA9QQkZJVNI9weSHnu5qQSNl9dSt4xoZ3Uk02eQHx5iMDylILukTRMu
hUSkJD/zfxDSklKN7JlDoDh6Q41EHqBt13fRuG8Jf0qMAo6AqhKHT1RhiLjbPhmlfP0/qrPnAuKD
Zm7V3Fpm65elvdmORgtbcU5qC1hXP07SENIey6ZL+2EBolCj0otsIwvLAe8zwZf3r8uPz2YJymyX
wof8rIpa73zEce0ysymwwVlZlIi0rKAZxa8qmzUv9KAxQcQjdYh85I4FYVxtp1q7qYbvBuXJ+fec
W1PRxZG3sqXEKjRAKdlzkai3nbsXOgvI8RCVu1ve+45qMKUFG9UGtznd9LuXDTTeJsfIiwmAlLmx
DOCTZ1UE7JPSah7AGaSWndihiOayCPLuVBQHG9qaQEsSwbL6ElB6o67ZRCDLvesSE4O7lFz+Ezul
nGNgPc35dro1Y7wrdYqvr4T2mXxNCDWGAfcp1JQdO4eK6uah/PiWC2DLQUVRgf9xf1Cauw18gOU5
oF1ohdOK3LkyHKbSDa4eUXcbROF/L2nFvrwoSzQQjVOXwC3KLqLRtxMhnBZ0S/GqIs2jPfd2YjnN
IeBl5wz9NKLXT6t/AXXP22VTZk5aVgeveIQpX7H8T7H2J2EbXc3FppzbBTPZ7Oh1JJkkbcKWNKQ3
1eeSZH1FxPQ9WKpsAC4uxXRM8+ityFtgW6j8HuRcjZZZczg1WYHd0zB4/HR1VTG2tY79309dUJhI
SMkilD1m2RkLUVmeFDATSaVxL1t04Igi0Btn+VHLZ4xBIlZoUsZ7zth5f4iu0DYSS5X23GOXEEDZ
J7/35Ub4Ylk6sDlsfqwZ1iQfpZXEELaiVo2Qb2gAwIT5qBInaFwtkfA1Xb9ZcxkbFecyzGKRvf2J
Y6kOlPcEFqLS/AfZEUoiOzKT0qwEO8CxK1Ne0AlK8YJDH5+gU8IInlwLGm7KLy0G5+EpVxVwXPO2
ysvwDUruM5GjaFFnlz+3pf20M7DQvSz+R0JT/ExyR1OMTW3g21ibFV3cTJ6SFZj2/T50ODkZnQ/4
X0iPvQrRLs+5ts9IdZ116bQ/AQhHFf02/xrjklqWRyJJp4uxK3Y0nX2dl1uY32M4YMkwqlcchOI0
Yzqr8FUh0aSViNEWDz+gz4iKSxRziKmfeYRbAgVkgjybYD3TI67lSgQk22Zb39+2I+i9/BSUeXxQ
wTyH2yUX8NmBIwoOokYHxYITrv7/D2QLShQ5DE0NQAf3I/OvYfgUuoyTjRJukYUWNSbZCZNa2eoZ
XdE/BSYr4vIkyt0LW7lNq2aa/ie7uDuu3+l3L30VPyi14bh1MfXSQhMbXv66UjN0bPNw33HS5te5
tZLfdluYmZNmESg+NkHnmuRotpPvRC9rUNvt1p1dNZzbX15MgF6lcucwaekfNo7lRXNFXGOkGRa9
e8FCDeuKS23j1mtDTBlZEhlqL87ZkK1/041EVkYn3MRUTIsaKy31lK7K2larzYmscNfbBQQPrpfz
bel08k95e9JmRaeUldLEQpf5d1KwMuM2x+Ofhcqs6CJGcYos9u3LZuJnt+7bfAfLXmXHVM+C7Ijf
Ok0txxaLN+hMUW/0iXik7CiodVO8kIJcMTAO2+ql/0H41oy+Km1xc3t2wmwgt3YEJmrqs/EKG+TU
f8vVOsicIBHok7U/sc2yjc1y8qKGcK+v5opQYNtoOlWLxh2obbywsbueCEsBaeVINwYoCynyv0HA
fSFG7nILK3MchOLi/n1i+4gjMM8fgpdw9CoVFT8ia7lGNkX0hHs7fm1iA+CfFIv+nRikOqNMP9gV
SFGgYS+hsubYp5BQgjHpHJ7f/IILhfBgt0v7sXswubO1TOunnwSEsHDNbYZqua6H59igSJTSu6WQ
B53cs08Ab8EQZbPCU+xjL5Djr8MGzWtiyv4URzdQxNUG58ScqK8APj/valBaUBNpcvarSePt2YoE
4lVPUDI7Nv6a5xdLp34Kws8IYI8LokdoexWdqmhlJNzkgBoEyiiBGQWQD1Ghky6GGF+Ucic9BpaL
nJzP9WTOUGYwVuKVP3aNGbg75PyYZAWvNI7Y6rj+RlSamxa/zaYZV0lED4ppgPJ0x3bNMp8j9fbk
+8n6P3ojyZx6grUun9HnMT4M3lAyI0r6KiMfO15GQHa0ldnTLy5+1uu4AP8ERkJdksv9csROsGlV
CHWdswuQvXDOuZVIsYrSqbLdXUnSudLRpAmlJvsM6piBR0QFRu7mhPS3s6/7x93cD/S5vSuLI0Pn
nTmvB9dVAr/XSldLgqq9zY/3TxKr/jNFt8ZrKLQz6BQqZ7hDYE9bCWM3J/ZTuFfGuX3pKZ9800px
QWITfjQ2rnfM4rod5t4zma+4597YxQuZGNWVhp35FnfRruxw8rOyH7b9lQ6RD8NAqQL5af+i2h59
F0iDthMkG2l8tqS0vum3hFjSC+MfadlxjsU0nf41xopPahTGA12z84aS0PfVHPLp1wn966+1La0D
DtRO4CqoYluCSBpgIKXvYvG22bV6Jutx7O/tCwc+RkJFTGuvJgAc83CJhByEH75fqGdJQBOA/5A+
4ndvNAuNatNVfJ+FjUbno3zqtoK1pEHo709rqvOe6hcQ4cD+6424smp3W2eoM+Ah9wpbO0q8ZXwC
85eJepwHpW6+rmcygQRYQ9ke9atCsmQlFkfCpDwyBJwk1h9+H9Q2JrgvuzZ83+bNOobY4NKUoXpp
wdgM5+GdeVHLmstSNuJxankFIlu0+Qo3zFFONg6t0RPKQ6O3IhrDS/5vTyKa+pVhauXA6c7PJFGB
XQc7/IvEYI0VPC2rGYe9D7bGAhD3LV0s74vBnN9btjhWBjw96UfzFdXiU+1Rk7JB51Jj9gq1Wfz4
rCwMWbnlc8rp31UEutRvTk5F6Y0CKyphbdPy0Ant9eAbBT6CfOlliS973dvj1VCJwHOkdVIV+LrZ
jroETF3r428XpX9IOifEwCaowp4p21rhcXIkcrOcke0eeNHO4BECE3K8+huODB/OYQrDI/E991Hi
br8mHs2ly2fcmsuCnPPQHmL3qRwUmg9/Q7MTEUNIlhfLtfSQbCy3HMNLHKjvrPsX+rM3aYr+uXAU
RB1SqODKK3kBdEA8z97XD1cxiH0b+SpqGSZjU03N+IGoXEv6k4NElYIhGM1lFPk78EXfp3/8Gglv
ikodG27f2h+2VkcJnpMcbrgalOfizLpnY0OcxNCJYtEey5x6N9Mm+D6VRfdp/wxy8+iRdEJ9JdYQ
HL7V3bjqS551Vmt45hciEJNkVNPNCVHSwKYpm3tLXoR8ufdlOClqgpPipfIqnPY0EJM6on4ROPgX
lW/YpId+dUwNr4AB6MHkVGvE3o+EFMQjBwvKpPcMvjoDG6FPThEe5hL2C5N8O/+9tTlUlpHX+Kcv
gIuMjdE/tCJqOmXiBqkZ7ka34lOfUrGafT3DJr8YR0vhqoDFpDXwfkr5B7dLFDxT2qEMcHjy3Ope
4ys4+NndM96kaJsnOmJahVcWupQP7lkdjnNjNzLBRcYRaZlyflZUTE+3X1IOCT9FmciB2xsM2hJc
g9O4pgFjLBoBwpdBTfNPVBPnMB/yCYFZQuTEhBNAh45ntpKor2aI7ZelinrSPvjeon0xlFmnhC5G
zarI8+dpLXgasviq8gxocGCbf/gh1lD5ju6dROSXggmH9KQlebocsR1VObq4fOOFCGfIKg6FdVMv
9sCzGISKti92873xniLZ8if3dn4AAMAodnEIrM3xEO0nkFh0rDyN+2usYfwl0KeauQr4t/Ad48Ir
Jq0EH3G4/D1TwVLXgGLCh/lQoAt59TAJOQtHy9aE9ERq0XHZlJ1Ap6n3BGWxVh+NUJKXhfy3q/Vo
GV4ij8aI9c/C1KP7VlhK+bZz7zjKJuol9AsIwlRwYGyCLdF0ucKUjqsb0Yd2TlTR30tXacbF/2tU
U0KPup+oBUn1CceKS1Tg/Rf+X24C3gGXN+9bss+nUtkizUduwPxCarURZwERYjAxiQEM8I1CakYR
jPEUi/xZvYPmscKGu/IQpRqcHBTEhow7kNcwOumftp20SUCE5nxZ+drCr8mxrRggg/Ld3A5cWqX8
kvmAb4simOLzpMolupCboKk3rDQoGQG1lnhPk3IV+2hD2DFJl8lpO8lUQDkRV3SjUFLBLPKlQdNf
cdWtBtW9WFvXbA4KqhNV/c3rruXbhHmmrBLG9vin+KWx1H0jvDlMiW/y1/2/ZXr1wV9CrTkhAN5N
JTJvTNkXAwVD25N2DuXrtY2ipByimWNJhk//x6yIIL1ECtYPODZH6oeukIEA7OW1k/5KIQ+HBETh
SeZQoBowVv/AtVBo7pYw1N0r6UsdeOz/AEoggVCxt2cfDnFtUzJ4LUfW76CckEsUC7Lh0tnh6pJ7
u2j6dk4OWmkMVQQP1MpWjZ8HOMbZRsHa3eY1wi9A1M+CqLWKjUPOSwYc9Zvy50wbHomi/pumZZ/+
oz1rQq66xjIL5qdUeYGmam1abjzt0s2xCM3aBr35fJCWwEZsEKAJge/fhDjPNVv/g5CCx5aOtJOe
eGLId21pqYAqPZ4jgaY1PUHiRQdVZmlJLY+KZ+A+RUIozouqOr99VubXTJlwen7OKeZFRNgOHuI2
66rPuxv9jGWGh4tde5ikC78q5q6vgOnhZdru8aHr5QDe0CmwLSV2+zLPXmdIXT8Pp0xM4IL/6u1W
N3nPdxKMvlhgcqwSf+4yPU/NiW6kC5G4ZDPnctz0kyfjsI3WW4MndtXxkczdsGCnlOSGjh+RZMua
R39bnTTbexT37+6Ut7LxsBVHoTS1DJop1xTSeAO8D6YNF/WZEgiWsU9EqcGLPNbyRBsXLzrBc6RL
Wig1dNJsR9/MzWzFECKNsOqPWPnxk9yvjQQMH7TtjzqWO3Sq75wXouSk4r3WOhLbcu+5qMZ7hifa
/WMRLh+x4rudnonQLv0kCNRB5smYD7fuDW19XkuB/vn39gkO82N/PtykVsDPUsD0akCxMnpcrVJq
YPdqKo1MC1BeL7B2MZ4fjBCRqLLvFBeQxJ7TPX0CHH+h831xLNmRo1IZqb2s4YMuLL3ddt6fFbi8
g290gNeJVxUtz4wxfKqGwiAIH0MapGHy9yxSxg5iMJHtww63gmO0Rqcl8I+ocpiuM8kEC7J+DApp
qiobAVhPLrO/w2JA5u4FMjQB23yXoPDaL63DQsqxu/WKfAZ69oDyXyQYFJIZMPdZXzKCg7lCSr20
iLskgSl/TQHn/jPXW/i/wigJlL18pspn5W4jUWgv94+WyJpn+1nAJMvHGrb4dQ3QjNQF6ZTI5PT+
C0c/HbkpbZBU+kFyTIk2/qwSf0eYlhdU25L9zDn6F2iCjVUtH/nDR1scXrgo3vZxkZaqHKCbM+g8
BPipPE5iT1S9AAK2BeI/R/zwsC7Uk2w15KQdiMzjXmdayO9EO5qx+gSyyti8Uoggr5sYjCgo7Dv8
hUCR/NM+zi4ykNep6bvpt0UILNZ3md/LIO0jC77tR7z4oHrLrOh4f56TZtmO5AUb+mmDYZP4PqU3
/fvT7SNtl5teH//gkbrwtSvN1xWMfj6lF2NZIzdw3pzhBi6l5O+NVH9P34tzC/ja2ysEo5DRSEYS
GNDVV9eiA/i7PQNGtRlHxesmEXWwc1pmvHKo27JWNpNl6GOlNngGh3xmYs/7KHL7+pW7lP1GzJrV
7w8/59I6e+c1RmSTuYz5U1jiMqVf1zRmrxiR8/LrmdzXchxSov7p8lrjXPd6+lHceeU2h/d/Rl8B
LQLv/9aGIu48oFXHFhdNUgkGs2B2VIPMwznAauC6uC7Gwxioi2cUfM3781W9TEBatRPyk855uk2Y
Kkr5zbRTmrhAVOZKsK3WM+cr08Wd40SMqR/QW6MTW2XXihKAflQ26ZLMlard2JoL+pVwz1SqMJT0
awnraRL8MeHPnw+sKKJxJA9ezgG34cqhlSB/aVMkCNhVvLSO+9UAvnaGfuXg6M0sMN7DUfqJhE/S
3yJlRVVzF9i3RyuJ3IeGHK3UR34siL5JVLiIeM1PEKV7XZn7fUfIA5cS/u7wA4IopzbFS1rTt6dn
7+zp1tds4do+jwRb7ohcEhrQeENHdgUJsLpxqYzhDRYpmOJuuaoDvZf4cAkOh2zX7Ua5E0HzlhnW
MTa9fNrq3uTbTYoukOUCQ7ZUAQpbKki73S56FtN5osU20/Vib7sPyj35R841Q21F0DSR2rmmwAvi
2aEaIoEs3hIILERn+/YMcO3rjukQUyDzYmF4kSOvS5IF0Qa3j2EEyh0B8qNBF3y8qO+DGnkrxQaP
ytabb2cmiy94BmV0oYMJ1BiFPY+85HfLhVUHYAodyefu/Zm/uoDYxxnvj3CkiQFp0OvCEQP2FjmT
5nG7UYrS++CGWq+RGstgQkUnNJ+RmWRqABymYM1GNNP4a0LhF9MFqMr+vmu2lWSgPyKyEYz9VaBg
dQZYiXYXPPBWraEqWz3QLdtqdO3NxH/c3tWLU00OxB77TdzbzbRu0uHnzT5Vvjv0FRFLXXJxXRGM
BTJdlMhf70JIyRpk1v7ie/K+Jc5fViD7wCEI3CwUq9O7Hvh6McFuPNH9L5N1mDejAbeotAu2fRb7
JKMEp1OSEvaU55SJB1TctB5tjZI7YGZIdnXXwzCz3o1g2Fo/2EY4lYjjA/SEgK5SPP5ssuC3Qtli
R1IbcBQCZUU7YZJaW6i6cpQ+lLtNfRY1tsPAIDjyAAjdNCEumzvyGLIrbCKP+N6pYZY6jO4PoFJH
0fg6mrQXO+I9Zb+395C0BYrwA4Gf/ZqY0nAAzUYKaHQFd1a2jefTzLvoLYwS0U82hc5AIa+DjHA9
+WuM3/DOoSsjKeZn1VzYGuzfFNSdhuYlpob3kRMPoof6jMxrJbxMDpDBiMEE7eTyQbCqeflV0OK3
G/PTrDorRc5NXg7Xfbtq7Du9/Pjv8R2z7LBXCFeNF2uqAMZ9kK0toLmV38pT04vujbSEqwhPbFHw
pl48gnsonMUzvoh8icpcHXC8nouTnsuLG2bm2gpVYt5OsANLjgM7LNdNKjRDVK0dr//GqXpCvx+/
T9JYPnmDpqnsLfx7vXLK0kVwmklI8WmEc2VfGpj5aoZAmRCsQ4hll4O+/Wrvrziajl9uFDRGzdtd
YMyQfPtu0sPMZcyLVc19CyptTcKGZwSdQxx3RpytX9FF9duoB1oC4oIqv4nrDiSV1le9HLKc9sX0
tAvOCWHJLkkryoZytVc1CEdAw0OuT9sy/YO/bAf1mooM0jRUxGyxYo0z9AmHy+7WhlF1dI0pg2oH
y8V8ruhvZY6OHPV+IkmktJ51I41ZxipL8NNOnYf9eSeBZPvCZ8cJ43uln+B7PAYK29nwdAgO+Ddw
knfsaugF75zu/CgoU9wGqooW3a3A0in/WqpLMosIGe5d6T/Rgn2eEJY9M4dQsBjApFLsKjXZsPdk
IdJhry8nYwVB1Gvcx332wJT79o4enML7QlySHCUBqgFWzoq+F1FU6dkwDcWfEy34vhwUzfaA/e69
d6DZQ7nF0EYQwHVEGYAkjnnwMYRHgvweKtlax+Q8XlsS69LD7ePsTlIslf+naVbL0Jo88OkVqW6f
KZcLBDNFlkCi79INhWO1yvAIiw0n8KCntLGI8x1UDvTqS0iLzbnlJHd7yJ99cwMapcCqV+6hjVWy
yaD65XVx+gTQVaAfngg4fjMBFaAMWmAOmxMZF5EV/nNGhmgHw8+O+Mf2Nekws1TUWTBBgUSLat5H
K9ThjkcHoysIc3aUtFjrmTULawpwvkTlVtmRkqtvbM0GeMHqeWTinjI58/4UQk2MkPCtzRrSwpfm
nJftTJyxK3uCdJLfZsJf2q2cY2aCHJvnq7JmOMlx/3XG6V+3YDeo9xaOt7XV6qOZ48FGFsbmru1o
ULl6+j3tRWRT5Jolo7fSoy1ifUai2FpGg6GJXJy2DpbSTpzqP7ZJYGBFx8/ywDKalMryQCWPcQ2s
iLl6Dfu6w3HxrHnGuBFor+LkF3gMtFU9VoL06no2tFZGbSj2llEbXzy921rwrn+vxXtA4pAIjbEU
acz3E0/8tAPbRtegxpm8MPmJNeT6JTu6hBmgYCljMNLSDkyfB9UQnQ5ZsLZFiR7AwIloPeJupQb1
emh2FnG1jzTB+QkslbJilxNZkgZfvtk9tlyxA3L9vNXq5QT0GOXQwwzTDtz2Pb6A6qoX2s05QwCz
akxOc2oEskFxRQsYZmYpQWK5Z6CCzqSj6Rdseaudtn2zZNTUq0CQWysJzTjc28op0uyKQtCOVpKB
4j1E4uQzh9U14/c7qHPJsTyIKTGhm5btp5lW8cjmTTk0al7EMEkaKJelCiuMRnbNAf48hJRv/o/F
kVFjsr4sanesXA1L47mf8EEouc/mCTOrWL4vcu7ACce44R4Dt18XMpw/CZmKsvRflZgEeq4s7PgW
kavFokXU8FqP9CFSCmDVtx0Fb64Ww9cvtabMMOz/7EHfjkipPDfJqlEjtJBISUdLBxFMPkg5cfRj
TQdWDuBGQ1i571BswWCluLV1fbjSWDJJ/nF71cjJk0/kcwZD0mn0fZmSsf4dib6pcubZFaAIlArx
V2gHtSsq2/jds1PqWfBrmL/5gUzVUJKlGDVC6tug0niXvLDO0MHQkpcNvQdZ3ur3jUIlJ2gLN0bo
wLi5/X1kzF0YJuWUsPvNl7kV28dOaSubNwra3E759oo9r3V7PLJwwkwGpVasF/8LvyT4dyJL5E6M
8yjhnjd8OUuo4YGrWcYfCbIq+uXBmuMgOdFADc0cN0hH+5TZxQlJDAebAwsf5/VkmQS0XCNvH68D
hPfAVaTbHqZ6P8PudyACjqF9S5LUnFkx7vQriMu9eCfgFsQe/7SRg3V6QtlP5EgW7BPq0NRyPsFv
ni+7U31INg+nhi01TeU4mMuIntwQac34GdK8iRYRWsR8nrjwhNSpTISh326Jt2P0+g254FNCAa5H
8j+6jm3clNDUgyCHb7hKfb5VLa1Jf3ACb5lQCMXMAXxEtcPc9zL6Xn6rGsxK2ODGe10gFW2t8eYa
uE/Yc0cCuIrgp8quX53zPLzacZYBQEymayPBT7Dy9g2e0Vn6Ww6nFtzaSpQyEbkRrqA7yI7IxpWk
ucPiRvNhLNZGSoTw95ATsZSiGXXGRHlI/zVKhjVOaVKgfdujDzHUu0QYZi+RqUYlNcBujaaOGT0d
Es3kl0HaeLL+ZFIIOBK0aPHGtbAdcqv2J1LyUn20ebClkJiQD3fp8yYXZQKv78P4SAGq8oqqyoiM
U0of94feg0OAClulECxAwOpKQJYhWvxQ1Lxi2tLRZTNvL5Pq1TBzw1N3Jya+u0diKa0fGchOx3Zk
ivhHOwPQJHI0LpvGodd/E3jEcg/D2wr6vgt8rINgwL87vrWZSRgg8E4SkfYx5uAaIUKiEEXBtTwR
cOqi8rE1+RptduXspzEjwKbfXs79qw5nz0GeSGfHCBju53WBm4PAHH4i09gJHmFQ3gQEOfG/9xVk
cBxnYG7SRa88pWelIZWf4nRSaTfub7qyaCgLYecwwixo8F6lrsilaYn4ELLpD5gTbdjVUKsY9nqY
2CrQnj+hOEDoW5yM5vmPhZ1OCaqvfme05Acnuc0ZyHH+2nNMfoFBpNUzisOojhbh8knQMgNHSktS
PcFdeajJarxlJDM7VG8+8V48ty2GS6OwXJSoHXbPg6Jl8mxww5EzYE3xFEARJYvmIUUP6hqR8tKA
UaYD/B2lMJofHz7erCWR05F4Uf3fF1+6uqDKMdZuG4d1HyQYAQC9E/cTqwSv9QvyoedsEA97mPkf
J5qYUKL49YbRWCgV9e7TgDG3ZdjVycErad95lX1gIYEuZ181wGi/PCjXLRYCHYRGfwWPGpVfL7Rz
DZuYMEX1EGOMtaWSWVANKV0QoVplWHTm1UE8a86QcC4+RyZPtNr8Wxb0rlX8FWeeVjVBPatE/z3L
BJzTSfZ2d5hYHLvpzGQPvzhezrGMZY19L8CApZueeoSz2NJUR7+gqPt20W4OppSfcjiA6UTjpN+7
YPzykQoGI74eGNGQlQj88nWNhmCtrJUy+qyKOCgu9dAMgIcbcKZIpmO52zYda6a2NkiQ19ajMAis
+R9YtyP41+M4dFXVmIZKsybrIuyIvBImUq/IHrTMJE++GUYe0LmJFcE9I/ipVUy9pb5VCaP2xkru
LED6aWAlmxYkBgR33fK7kOITs7slBn8PM6h2hfFvE8rAftN4EBwAIMbA0nAkPqxVeP/fPFnWZ0ZV
FNsmLWYAbn9eAHsLlvhgIQrdrl+KyMYJYCACmWKEATV8r2jWH5qZrzUfm8buFfADT3QNr6Wr2sfC
PV82kt27fLgLsTBywHnFccZtUB/TF57PJOETw5LjK+U423irKiozrDh3B7Fc+f2Oj8LSKWzqda/S
AEN3DaasayKehYRPcuKQyEdO4M4LHCGTFDs+lAaCImOcsHF8QOU1/dO8RqDwOnyx2phECC6nFpxY
UWJ+5zENOzMxb4fEjtle/UTAbH3ibCADqbCaI0uRG+EfdlEfaZrZkks4Zrcc5tckzy1HjfOBsr7Z
3it5E1NRW9/TDJc1GXWTlQZbujAqkOJS/9Jam8VNBVQ3lrMqGNFjrI8k9o05CwUmZH1Nn2snoqkf
LRCoYcQdujcwT+2xkiwcNT4BQ5uYrYiZHgUoCW0ngL+6NqiMNjXk72dJENgxIswrP1RAqNnHT4JN
3hRD3HkdSV/yLeuJpZXaCQyoi9dORvDZKSiim/gIVLFgsGXCnKqfwsJMPeo0eSKGeXQYSLc+LZ97
rwQ6qwHjwlOx5PN3oC9l9IC2kWRPOISEcDaUoe56mvT94x1nivKX7u9mJWjB1jy93Fi8JEY/hjR/
mmIPAODAAryJNHtEavLqlUreYreKZtaJBhhAWjJleZ0LPVDv+LI9/d0bR7dKD+KdfFKH/dxWJk3f
PvmFBGMQy7NRQXeqHLy8x+kRngyxHDZtb/sbkI26DBJHgWdGRksCt3U342Jti4EpOiX3JHtCc7Qc
aIq5ad6aOm7Bg82/smpBbfFoTks5qkZ7mPxdEOUWFnl6MCpvlBUIYjnBRdIT/HyH2CBXBXili+PD
4SHpAuyeOsTjI7V/veI80XnQxRm4cwSi7vjPOqYYwqe6K7QYj3tyaWB5aqxX/Z6YZ+6n+8KzpYry
TABY0qKuCRqz9xEGrjwgJ6oY3Ov4CSFNWcQWaHtmHgTnqhfSsl7RPV+UB0swzGRbXSUby4fTpjLp
y642Z/oqZg6drf5xbEUnX3ENQgutouYZaLTQFx1P8neb+Dr3s+U+4bjY+6q7xZDioxxZu4B+J39v
kF96MSqsZfdMxmNYiHnYWzp60MzGsJ2e3twkA4UDCIKXImWO6nMDouixbXs2/yLfAaq29nvb8TNW
zKlG4MSuTM+cKPVoJ7ZFjKkzmdqCLmucsOJo+pycGX8t+sDSMDRzHuHCkfGJ3NczSWeVh4R7TKJG
EVhRNUK1cwWQQKv4vSgaJcEzbvq0ZKB+2MLjnt/mI/bp3uzJFa1Mc1VzIcgveeR5DHtWX96gEVTk
GwWNKXesqUqeWsOi3MGU9JNw9GAL9maMhjc8g4KpcnFquuqaexFtIuddqJ+0J4l1N4XEeyEq11nM
Vi3IF45xFl8kG9gwParvm/TJg0A1Mep6RKak+OUtchinyUnW6UVT9vu2RBxZuzgcDZeas0/u5vn9
1/6R5fwsCS7j+RpeCBGBvagOaCAwOmYENr1Y5aR5FMIz2Ef80doYNbXoNok+tHQtdYtjqvGB0gwd
ltMdTOlTfIij9yhTlS3akh/VfN/xRqnr0CF8ffiDlbNCsLksrqgCHJzkf4sKZY1FwppovAX4E0d5
oo8trxJhrUusQnu1j7x1m4N8KwcuhDZNq92PlefU6FgRhZ2ON5MpuCEDiVk8hr76/+MJoEa1xg0W
PgCcO7SEI7ytFwfEgXhPDrn9eE56BB3U+WP2mtV0g2OeK8AOAeRR931CRYy0Dg2fPg1hxGwWIQ0Q
o+3FlLNREKlrBvsbXMMOkAB0/a4Y9OtsTWbizhfjf+/CM/0FsCdJl9sWSF84ZgvHMRv+fAaG+hcw
zkCMbaAdOHiK5vSmIIEDCZeNpUXpLDFVKjEj5atJwR4AXedUnt13EeAOHJxrIRVDo0Un/exZFvsn
Y8E/bMvwvW3wik3Ys6tZJLSwwPQ1q/DhfH6l0v9/PZD1W7qHV8tONttYY/TX/4LSiq38nXPirDF7
3nIFVI0aS69bQQ16o+E+TBYtq82j8o/LfO8LzLTniRUlmvL1fxEC8vns1s1Z8MONyiE9kZ8zyt8p
mnzqLbS8ygu909Guabai/0BIeCghIdBnZlZF+PYNfPRQ/Eiqr5aC5F1zPNtEARUR1YYmWHeO/OVL
Xm5G96uU4bpSq+wPIYRKtChyIZD7LXM3Tx8rlqa5XOg2pNnGw0aMTR3FPp2QZIu0vAiffxtQjVFe
o+yJmDmdue3zOnBJ0NffUxC7s0oqsGlVWo/VzEz+wIQL2NjQEKcII3iFxkvuR9CjKdxyuOx/7vHb
gnfaK5EHMRQqW1fX4wdxmELxm5yG/yPAM+NjkRrUZwSOOFkGHxwz8xONmWQnvIg+3kMgiFWdXMsO
XW7hMdFlhKbWz5Wt3QoLf6RsEdUGR350f8Q0n0HJlUiSZs+DkpRQ5wi3Z7BNmS4cLeoI2m8M9jvO
zwmjNl8i/6JVvd9KCstFYpkuaGWOYI5wGVtS8ekxnYyItFoUH2KxWsMi+3ST+dYgHmbWQ++W98UV
lrhu6pkw/8q16+iiPGwqpbE5Y4boJFyZLPGEAI7WAuCAbjRtF2djg8yWjziatPwzXnC8+LSB3iwR
C5FUxm2Z7KO2DXHR+y8HCKUfBolgBYhskM8sGGRsXx5SdzR42mF4SBqHauxXcV9w+bOpX3xK+z82
haU0x2G0YmG/n+LgwP91E/RLAQ+z4cWFx+pfQYyF4IbRqP83nFe2oEDqLdnkho1jZ+KWu2SjxdlP
6o+kan25BKpT18dVW3rO8Sv+miHGCmHH3LYoKzY/3OBllXW8Up2fD3orV7bsz/PLaVlD7fC/6loT
HAsxT19q2SQHZihlVZBOhePAKNOyoePDeLaWEw2f+y4kF54k17ewaq8U4aD8vOnhvj8ME39+oaqN
1uvL+6Agjg+0m0LVHYZAuUc6HJ7MgVpLuYRcUeazHuHOWlXrByqx3E+mpbEs02NLLMix69iFzjvt
vtk1TmxfLiokyBUt6SeEslZA5gsb/Dgs18NjKxg3COUvyyHG77HFskpHxdU1lpxkanHwuBwSmJ3J
kQ9e1DoT9zXg29CzAyAlRo6v9zpdKaZ9Q9VSTAKxDqzU8orlRD6BVKMtUjhjdkqH8fpKHauMlAiG
SU4jgo/6UWzfEPtAxyQUyl5QXqW4ipNptIWiZM7/g+TO2ie5Rtc8csPXOBEsA+VaIWwgfCzYGIjQ
UoIVJYKB187Pa8TV3wHtFk3ua3dym5n+vKdG/k1Y6nOQ4C0YEtbog7wH77UFr0d3aVRFTUDf1PCn
FjKckFBng6DwTIqRuc9qQBsZG342PO7JiyCCQBvze2Wzs817IdgZRgtD1zHHN8A6gVyKlgm8jhy0
tkmlovlw6SH7VI6uoOd75+jYWXHsiAb4dH2tBzcHiV4982uXlm4SuR72P4nO8ydRLEYInTPPvz0T
g7crWtiG8+XQF+L3s830Lvy2PPrXCweELHAJQn9ExU2meINrOt+64RXmJMfDK4Hv9TXDuBuurz3B
P4aWGskW9ERoXva62pQyxnVL9BjIU6ipFJHL8VsUcEwHW11qpRZP7aLUNroNULS/DaeL1fTRHQ6G
XJ3pmTi0cwlKzVqc5ga+4fCOARh3a6RahdC+PhoedMBoMpmXNCG0Bt8gu1Wg0emspfz+y1uImoOi
vw3gazNQtpBDXQJn3svXzm95ehsrcbVDTOU7RJcBlY0pSGmMMwZgK+B5k2l0vqJFo8HCGWb2wQa5
uxuPTrGUaGuUJlADjAC+PQFasgxiXFZW6eZSJrC39BERP5DihDCOhRyezPLQj/giNHtS8NQKNNsV
axcXC2Ph44YeFO/fvCT/bnA1EzjWUSnBdhC5W1ftHbJ3pxcjTu1IBNBbBrMTArlMQ1jLshKt3Cab
DDnqi43ytx3E4LBmbU3UOLB1wrSaGWjo29YUGIpt2ewUVUJWhgMLj8AASpU60pNp51ffTC6OF197
x8SNDLyTJ/6uUnZXx3r21ilG4y/1kHw3TIFGT8WRBG8m+G1uO5qKAtTBOBLyYys+mRmEC1ZibRFj
4sMwhIq050WErcEb4CnNU/RTWYK001pFNF+5B9vpyymNaMOqFZuZlixUP2tssJAAIMS9v1Vvnenh
zMZ/F/f7XyTurz8Ail48DrxGMzjyJeM1cyWdgd+d9eqANqPTvhAj/o3HPkgbI47Lk8J6kwIBbyoW
5IKB2+O1XGsi6kk0VknS2O8qmzC+I7Wunbgh9bnQ5KVtO0bQ45Ck5ILImPKmHI/MxdF5FzblER42
XeEefDLi8Ac4+iAJsIRPS0qdmRNGyjoBmPq4N947vH/T/nQaIcfUBF19ksxB5yHU8bD9xqpizcuo
RNrHtURdYytlispWN3CkgV/JxU1KgfVTusI8mWbWl+WEaVxB+ZEhYJvoUJ1gP2C/Ig4KlVqC+lF8
vm9iG741sobL7sGTrTc2XKcRnc+GObY3X879X5SuH1gQRVKQYmxCHD+f1wFMFpXBHtDeM6SEVbzV
FUJeXHNQACS0JMXhOYZVuSxl9zaXhfRqFzWIN8tBIepbX9JTaeTHnAXZwzLwW8mkmF6g3LLE+ovF
Z7CCOxnHxw1M4wojmxJS/kIOeaP6q73Cw7A5qflgwUSQrJfiSAuxWCGUtmOciWJCYVItCM4WW8jq
HGQPlhXTZtEa+41dJb51JeD2N2iROShTklPEDQccTaNLwmXxokoO5eqPz4ea+cIvoai24qNOxGXM
hRFcph0fYuBbKCSKPbk7Wu/V7byJMJqpeND2UTXlVGCTI2ervVgA/DY6WFsjkuoyV6tgVPMavsZH
IbUw9JGb0YLY2NFqaHl4NjCig89SNx3NPTukG2/Dm/v61ms5W5co6zRf7tZ/qBtMkHfgJ18MCcEo
hDT7FkBWBld+fZ3BzeDieAky7tMj6odTtZ18LVcgA3c+dFIrO1V0pt20mEZuA1oWxwsRCTfWkNWP
40j54N7ceYmD/Dp3fr+YQoGhi84n1df+aQmcOPmUbcGUo/f8TH6+iXRRyLXGKaXDJhh3D8ToRzpQ
CNakyaQuWWtdXWRTVemOUSwW1HkijTrdoqLAOrX5tUUuuzYAvpMzidKHtnlhGzMMZT0CZyayOBfS
Wd+aqkwZQjKAmAI1x6IYAhoYc9dnJ0pI4PSr1NybWAuWGwHbSY5A8stchSHPko83qmQK2qP6NxHe
eaeDB5vPxeOHFEj8q1GM33YrSBGREWA5XCdgoQyAky2HtLyuE++yEkjeOWzG1DSPifYz2Uz+dRtD
qpVugfl/OA+W+4ZQNj8VqSYeduwfMittTvj0Pari4f06RlcsD1TMMmoeh7RiWowkjKS9zPszL1Vu
OR0UNgDH+4FsCyLUIowAfrbPMi1jY9wTyEZV8/vQEGASAn0TUA6lVRGxp3QGY2sb6hjy1EZksohg
UgVtGuOW6o8SLcGy0gl3cPG9CQapPtjCbc0j7ajGj0be3mceYA7ox26YcM4mWC0VaaBgyKUa6pq/
7SRTjQn2yOK1rMRytQVzP6+TYM1aoi02TEK0FtlA89I40NI7+7v9ocjBEqsQzcmnzwimlb4wfo3Q
Ik2mfnd528+rDC1y0nMkIsxeMnp0ZbDuz8GOCdW4Ywy//FF66Ab5Bk8q5VF147FV30P20sUygsj4
W/dRDFxhyM7k7sEB0hwZiw/FLI+pEn84xTP75Fx4NTmBoDB8WmwRTuufxXIUrdFdO7DFzFLcS3or
xQwvlXF4zgwTzld963ml7u5De+Dmlf1tAzqemoYluAGW9rOQRJzKyZM+S6wkpr/bMTnjSj4aPyFr
O6PJRYiraJectSk/a+WM8RwMGGxvy1dhSyck0OmtblZze8xQYMypHYolkaCexnvx7MODk5FXoDy4
96ux3FA8Aaoet2BC2Uoji4imb3z7IYcYrAg4jP70vylyYaG0jQ/yjVT72y1v9gNZz6o3B19nOfzs
TpB5ZpuTxuRuOGmRjN+PMAzRcVaD9tBzvr1IRVbEtcrSVZQWL467d522maWOBOM73o/KtchuNUVW
qWj89eN17zhKbyzf8Y/m1ac4dj15w+6TuaCnrEpicLiIPiCreFFSF1+1TB9Z614SCH+J2kngdgVO
fB7jUNUbj12UoTawvnl6AyIBmmTpC7ouSN6/3F9/mHxeKZ3yFGUsqTnvl94RdC72xyv4mFHGl0LI
BC6jbRr85/YBdtIi+GpaYKdEJe2doczoEkS3Hhj8nl7+Osr7O6hSwJp45t+BanHZ4TEG4Yp0Nd7f
zoaCX9gxbhgpU6oLD2d90Ms3ukTPg6VG26uRPxNQXF4JRbiGYN/1Afd67Wt5vR7QUXMWYOo0j+FF
qSqa2pzAcXgFKz9X1Q0uuzREhIqjojXHWD5AbmhdeFf0+3OB5Vs+cTcJwrPZ6PoVNy7+cxLqu7AX
rOCJZG7QpdTzqucxqdxwgBI1HKDRoHZfIPxwlNGMdTLg9PekSMJNA55PK44iEVkucSBnj6U1w/Q5
V2Uf1h82FrpCvYzWGoi9Zu4ziA5Snz0Z9f6YRihwLqjXRtIt02IdvtoapBA7JEwgc3mc9vYt8kD2
FeouFwZkxcncdr78JhtbxI+kc/k0+17xNRbq3smG+f7nt1+F7CI0rxRwrd9JJmZAWC79bF8CVOdl
tARd7eIBKIlkqMjWaYLunmgVhg/AbIbFKT/FqfXKCl2M9zT5b0DUZop73LrExoTH36N36JMlPqYK
7WrPbTcZyWororu+jwgoukCx12GTUKmpttiaZbfIfdn0PiS0W2cTLfGcLljvrdBaFMzORor7dcc7
SCK2n7t0XQNrZDYsW9sYvUdKYX4ncaoz/rRMXuCKRwaYho+oKcgU94WBNXPjVfJWfayZXurUZBel
Ay1kWQT+Z9XDfWsq5ySy9+pNOuX3d0vOrn8r1c81Wf2R4MCmYAYQoAnyK9DIShNB3NIBmWZ+d/EE
Y9KrdAqt1b6oI4ZncsJbYkHHsx/tg5W3DpQpVVa9v+DbGNo7tPcYj/x/6pPS2aV4Eg7QxvQTOKur
Nrb/d6fVCMREyOD6GcJLmvMupaUP2gAMMM1q+wvqlG6xWMyG4lwI2uc1QkTM2JYgoCpE2QYTl1ng
iBuYjA0donh2aDB/2mLJwKGaSKq4HXpnh175Eea7270HsV7QEtiUJJFuwDEUwqZYPkwzh+v15jXp
bih340jV6M07BT7ktFcu1UfQw3/MXQ+MOAoNjwkfxnR8SelnFmbfgD/D9HRHGrVhC/8tmnMQSCYY
PYKdWwUcP6+LPt9GI4dsgipLevwyzAqE3SrOj2B7cDN/ZcopZADUn9C84PdBuC9OOb4tyOEZcRYt
PiKNl9QmIaq4dwAjwPG56x1xUXV734Pp5NQLHSpFrVRTWff88Hp1c15LWclHjZ+bW+mtxNDh8cX9
5oViM8pdZkhKq8l7DTPmeOelutw6DvIFY9+74hTZWDnF+3Pq/e+i7UEI3HydXqRdG9JZytcYx6/k
y7Ss1f79kmMu1EPKvf+jT738ox6VR7TdVRbofOpmc+2TTZboVAXKSl9nsVazwLgZQ1lV3D8lJqfK
nne4tmcq2W56s6YXG+BohUezLVVk6ONqz+gJIjtdcT4fIRU7OyHaIRtjFc9WVAqXDnsRbT/0JquZ
H1T2Fv2FEq569pHwLRx1kIzxCxlc3gaWSvi/iU3EQQBTKClfi2msQBnRQ3GUE4MMaWRDZ/nUnroE
VUIRwL4NR0DxSQjBe1A1FuDDO4G8ksPDtEcZ6gGb+VR8QOGY7OsfWWQictbRijIcT2ELeoQlEEqN
qhXnWf888ejBOEG7qgkwp5TkHIraDUBdaCSwmXXWKhX03ROii6Drh6fi5tdXxBifQGi4JTUQgdl1
DY8e2+ow6vEo3EbNA0AZfXO54Et9yLHbU2Z85dEduWGQUdGrPgrKvHf7Uhuk+DwzYJKvg3AdUfg7
fCxGJYUC0ZQDS9goowl+ndX5vg3wvu0zklx5WpbtldnghYUjLr6jfEp1Rcpv3yH6dNtdZG0sQIyp
O6sCPbfJ1+Z1NsFzD2N/vd2amy2Ojx9gYeJwmTxeCR7U2zPrplnql1lc3s4rTewNQhUWLLAn3LO8
i7tVKyONqzoJ27Ye3gMrQtw/+LxMouAr0HpgA0IC797VEPKv0mzG30fkVl6CSFWZ9p7FPv6wSJMR
rpRfpiIttmtMHAhVkQ+k96F69DDVFws37GFVQwTBvX4VVVoNwQSEl2b+yvb7/JDfI4lSoNGsa1hC
ldyE197WZRiQXNbEnKpTSo5vwqAc5QUfYr+8Vavrz87ChNRg7aY/c0+HtY5x6+psWQbLhmftouHb
eR6gaIpHWXIlvFSERkS52frzBCp2Y53S+8n4qHIbA7ZCLITNvLYj/MbTRuLKDYVdtmXiiazdpeXY
4ZVtdDa4SEF1KMKVYQCb8pWrKJrrR1cYw2MkSMg44ym6ydT5/rZ2SzMXQRTY+wDbszBw8zq5Stjc
8NNETbV+XilrAhTmay9upWZ7egBwTzsl5U1aKqyunqCuhdsbNgTLzqYTygZi58C4XwVQmFnTg1GV
xKs1T7/gfBJXPzUie+S21KIIpGxp7D3wz1ToBYA7OUrvu9QxvRR04S6MF2CQ6NeelO1sBccPTCNw
jQvQeZ7W4/ZfpMxM/QsqgXARBKn0fJiY6F+tvj+VJPsm5NYkeiepdk1B1hl4zkc1cQq70+2kU4cz
DN2QyrNMkqQO3ualPVrPsgg/A2ndB/s3aqqzIt0dHXkyRjhwtN2ihNyJA+r4bDfXk8+kGvmSloub
0V13LxHNAmyCSRJ6VcbCaMtqwyUl018FjDMusGhOuSr+LfaQJ9G39YQDN+TMyasZwPZ/3oKDBZbu
AHt1VAJ9WgsSdIJ7JRsQA4wqRFIQV5DmlUlqMo3HZ2ZzPo8FYWCchRoobWKLwtbJF5eX1IBBwcLP
OU9LVEwoOKD6WKN2ltPXEJeGnR8T3lMX06YdcPBCKehvBa+wlgmtKFKyhk7Oe9FAyF/Pw8MnNwTN
wmrNQ/TfKgPcANFnEce4KxudDYI+B9uZqLCTHMgYQMJiK4PzygEnEiHfsEBqlzuWAJO0sKFrG3gE
7B+icCsV0CkyEU127KXcgl6B582aNnpZxOz4BqMuAOdiH/InGrx1XF2z+GVLEupLLsy0yW6jMJXo
NrcfZ8882nM0fQ5RoMQXHu3lGC9oTnN0PPyOlM4v+BdW2AYFqywWVIbKiD7/xHwGguqP4PPlMbiN
AMkUM/RJ+A86YUifRL/0PyAiEMsQAXdTOjvAd/lxo+v4GO6tHL+NfxyfW2fBZvyEq0KWZ2IiNacm
/z6K4wTNKFH5NII0uEKOD6/nbaa9L4bH+4+iH/pH/EzDfJv4TILZpnH0uDvbtOMQxeibIXcUk8vH
y/7Qki79bzdXdt23CxvVKlSazC8YhxDHPttMgihsiwvbp67wbFceK0bdcXikJ4wQPR0ROcGt9F+3
9NVj/39FaHtT9Ogz/gWvlxQRnuxAhrQyCRzd1Zy9gXpofsRI2oMtD5ANiMT0mtmh9sVDVWITRMq0
pQ7yqABpJq1XpM5W8LABXEPEX8m1xYaUMpLNdTtGuWAnybx9NWbaT/AtbTOUjlL7Xem5O4KydPAX
aIV9MUI+AWFqQfvt5cjAPCdM7nflHHazK9EHP3I47V6At97Hkwmn3Z1bHyAuLJ8m7BqEcj/A8EMz
igrqTUAVbi2w5PHfI3eOD4Yq/yLsauXYmBldJwmAhVMNOOKXzITLb16d4psFrD9IhyvC6ygt3fOJ
9agEq/9k79ssq56EWF2I+/C9Tz9ITyb7KvIL4bEr01w7pXOfhWxH/wuDNOyxs7dux+DCYzIMMRwi
bJAEHkJ0IZOYm7fGpwAMvHxlH37uPuNX/sdg2Y6O49VdhEigQ+MYOOKbDE2lhtY+4V3WZtjXWTU8
ck2OAbPbJrwpjbMLvzbYieFHRZPOvtLrDdBnSlxKuSFXkuMcUScpfOFuBnR5QWHtbVDD1knTt+c/
gQcEpdSIKlvQHxT2ub8aDsfj2s3Euhu9v585kWqtc3S+cTdZIfaItb3iRPEOgoZsMadAoGS/stMb
6xRuDqLGQaJd23q1WUQ+p/noWQKTkn7Jq+Ggu2S3SL3G4G70r67/TBIFowPgOR8tw+za/BySwlnG
E/hHGdVoRX5P5TOEVF5AyJdorNqbFJXwuIL6gRBk5PJGkvxzA6qsU0VdGY9OBN4Vbj42FKa4Nedb
taIrF7+/iob3mxQFy9IwvNJoHkIgBX0qc6OZEixQnCbWFVLLv2DHdsQj5s+RWTIY3ga4s7levK7g
/MlrWy1C6W28je+oLcsq9bNPnt+Efm7Z4GdnkNaE5ytn4Oqu+QVrWulwgfUVQFbLX9COMoyu/l+r
p5tJ+H6Ekg096j2fGKLohQvE3w/mFWQ0ncGaIO4rgaXcr+69Th0VDdzUzfVjuCNoecew4Q/dzJyD
vXkm0/i3AJpT3UwekBRthqAIWkYjE9jZVx+4yMoAtzUR4o1PPcgUwBPPGcCeKQKXqOtgyklJsadH
tsGHfhaa+o/J/ZlBpJmJOozQm7Y76lTLHJl45rDCFkD3qFCtcipiADL8H1riu8sfSssn4np5rZ6h
hzKrjdYmXeq+dc7aLqMMzUb7wW+jAIRA2TsdsQlMNfXsE+A9cPocn0+WukrBoPl7ZmrmAVU9KsYA
fkOkd5h5BXRvLzlPlnIJ+Pe7L6Cdfm7S6rhnun2FOy0kGj9beQSDYebODGtAAF0jlIIeRxG/WiEL
gNG8cyCiZyvmgQz5daRd2IEVh2YwNfpeBjJqq82wOq+e9TbsWcX9Z3Wc3KjVRBDockHgeoZaoyVN
h/wFKH8X4JrE53I6cpNh4pJhv9OucFgZTVzWcvn3YYwXzV8MOybVlorAx9IzQvy9mnkUNEoKaRna
62X52BgfqqPtRw2RcqG1hdE41gBogIMsSRiZUZFVJi08flXhqHljj3jbvvFgfkUaQKiLsiiRcKBc
8GJXfGORqiGYneIhizLSeDiKiz8kQ81ezlplDUNpuSOgcQSQvu53YYWOO5DPOhY7SLUzlW6i7oE/
YDlabHd0Af64jR30LR+J19OnybMyaZVfFE3Z93COFoxv97wDaXOx0dDRJKPzVkLsI3KrsT2sKbuZ
/0urb1I0bpiMSa5pO28oQnsVLxW5zmYMec7sij+SiqrhTkOQ5SRdBvmfw3M1a8kL0PpyUhmGn081
hMgDe7B1dx/lTrVDZ40PWoxTZhxXzwrURnfONWU6Uc+Nr/edL7ypnp8dE5vVzW4d4dNtETrb6RFD
XbaNKweblUG06+IB0DW9eQEC6gGQtu43BK86nnpiV8xUOk9K7AFAOirSZ3/8n1rE9K942OrM2lMS
WQ9HUWNHljNDJvH9cjgq5M+HRY4R75CKlcNCZcY4SV+YCCLp60sZkl3tzVWeOHFy8lwhrUqseHag
QoIOYfPXrvZKUyjZT+cmDexMokR944RETmUPd4CTvgWwFe7vKLbp5EipnJXOYnD2YyZ/Pqq+S5Bc
7/Faia/Hz3LZWldFSaWGZVk7DG2pcLERS/0p8c42/O7HzH7Gfj+51fkh2mdc7YcfGBAYAhNEeNI2
Zj+dREcdAEqSukZAElguZbsftiYS9u/pXIaxyY6ZAf++W3FI5CN65hHR+TZJJO8JjX2yUG1fnkHE
zd4LUhNr8J/S0a5UY7B5BCSp2L4uHdkLg+k163weGpw3fWgeD6F109MAr8C+E/nvA9hbrX82QXPF
Mp19LOlHlvFVkNJ71RfGybgn8lkqRv5sGbT782ENHdbvOSP5AXR6cI1jHmNCZNw8lrgzclaRCnpD
vvZu9MqPjFpjxolrKjUHwB2whulYgIvKYW895g4iwLbYGtVX+YfzRrDIzcLfOGXJNl2S9iifxjab
P5iOtd5gdjZBdgFINMWlrtzp/Im9GvY4rDjA5VuR3ErHzeNozOvF7LZPmGtBGulN1WKxZwprurMo
fES9/odasujnaM5w3OZMoxeiGYVxRkfoTc/Q8rTBgdvpDnPYuC+uPXzkphRYKYYtn1fkbrLE/Uro
3r+Ex2GXnsOM4cjRcmz+TtzqkaYUAFe4o+LMXdUYRHgD9dN3ON7BnZvyN8+q1kTlR8aX9b8oCEUV
AZalFOW2BsPHh75O/i9E1/KEXG3ogMli+QDxXiM6uvYWsL9O01rFKu2i9thGgTv/+uzgGqFRWyGr
sNh7EUlFgHzoeyZB9aiE4l60aHJIqxeXl+uE8BdDj9PPObWVj+fTsQAP5QfTafFlQZyJKEw4rE9W
XlTmUePFPRirSfPVs1ec9ndM5b27eFoi0L/SWdfmSePlIyPcqKDsLjOgr/vYbI6eRU0Mg+9qCYEB
qL8SATjL6XdxWSj7dlihRUyzjCcUcIhFv7d/LgrNHsglQNcdH9mpIEO5UAUbviNa97eI9l0SAMgG
aby/2iryF1a319q/b9z7tX84rdh+oMY+X09nHFF3QozKa5aE/Qtlqqdx1k9GyPh/o7UudvwkCuVc
NNx4/qcPYVvxUsEdBiNDhbSRoAp8F0+xqjQqcc62Zz6u1HGgVXLervWb/RkyMPZRZhOfM7RQUZw8
vUNJqPWDBiiyXXLzo7D+upIRKrCO4qk4FaLwEt4RZehsBsVZgzk53secEshtf3nLO4qppcdmELKB
jkmDxtki8HZDOQdwNEaHpgK8AC+WOH5/HV4C30NAdcJpCukUzAeq77ygz+y4YFUK/UudNnvG5R9F
/2gqgMXkMjNuhlscvw/Mc/6QzjZg4RD5k1t/d9y0vg0oDDJjcNUnLFhukC56jCmpYOx6sZIcjXWQ
IbawU0zT4LfsaJuWF269UHbSmqy7LB653RaRIb/l01mLrJ+fFsb8svhTY48kas8nZXRkD4nReBNE
uQZhQ/Ce9BL5+wmsWptFnxIU9p5OHWzBsYJFgsE54i78TxwNERr3mWYvUKwXRyNg1b5T2oNokEks
7qVHChykyr0ocmH8G49AwA/isWn6BGzuYsy0VBadRhDbsfB1hdLj3HQa8ArxScvYyZkEhNRAbttc
lZgfN8vo1U90ROh5+ouUnEpaLIqIcfFajqT/lsUia5O/+itBXLXHYZSs046abJ/H5GBVhlfXCnVo
HOR0BHFLN+hik2NsKXWsazbCEdQGg5BdHVFP3xYZd3Vn4vWI3WSrSd2Ssd77INkKzoaM8YdBuCbf
G1hhGS7msbtnqiQv8L4B5f72ifoXX90Dhe6ley1HN69aBKXKDllBMTxudhDHEi8bO1EMjLwOorTA
4hzqy0ZnFBjzOwf+qe3BHepMUD0pOum7hXJhTQhb1c+iSNzp9bK3Kmkz8fRUgAo15mLOHp0hduHR
yMIF6l/PDPcuPFozusmsJx3dgVStBpDHkrGc5T3bFbhymGhB3a4qXXJEQ4JYOJcExchjqnkjxjF8
IPmnC8ZYUq8AcxqcEPxNsWeNe5OI7NoAQ2Vp59JmXfrkVFt1koa8vH2EZNBorHRMjACY0+4e3vl2
GMhbSJPpcY80BTBds8FifdDSGhtJjN8WbYmy+NJEhxBG6Z1b4RiGQdLGgM8vtC3+RYNACr9f45Ao
jfhby7UxPn2VShKjbw4J6M2x5wtCIWlPecBkrGRBaWPL3EmeXvmdRbjT2LjTgG4CTqqtNIglAGZc
q2lHxuRa1LGGd79yGsNHdGruES19jghQD6EDnhZARHwn3gdwBVWJCuXnRrsUEU/kyGKIKEpSW4QZ
lhcdZKgqW9iD3SyVhnUKtc9pi17pDdo6u4JvCD0+B0Onu4B1zy1jSXcbMMad4HjOWxQA+vIrzsEP
ZwU5cUFgT4DXQcy2Iz/YG12/zAeVRxnHBs5zQ4zfxUooO3Irwa16HkmlQHzl5GgDyccWgG487IRt
tdJ3Fsl7lZNMSzqL2dR3kYLW3o+dVZ5iQcTFLm6VEDt68hNIzk3awnAgXZglJXbq/Jb2V2mIm6bi
OvOnVvvigzbll/ntlQbe2iDzOxLKpzzL1sLSaOCK44lQVHx0O8p9qEJ3Eb/XD607LHS9KR/lot+2
bSRzKrGfPQO+OeCX8o1PCNqAlmGoRJcMsSt1Fkkkj/fbMLkOptF0HfKtNT6BVFvcOr5niIfHQesk
DxqF5WhQgN3bLmXJ+tKfGsy2Fmj48KiFKqMdldVDJW2ZPjd6BIc2Ea8uSM49Zfk8qquYbWm6I1Rn
Eo6B7LF+WGMXm0EcikDQsrdNiJXCsXsX87f6fWP3eoNn19WhffYc/Nrzcq8WUcpolymzMbWGYbDK
DPP+ePQ7AY7u6IQD2dLzENb0q2fgmURslMZSQKlxu0pbocfwrtIRYdWVyWTZJZjQPWclFzj76WV5
TsPbra4o1zb2KhBjsGABML81m+CTGtAkPU7ErOW6i5qijCMJLui1HSosmw82nZxrYs7zShhS/WeV
/JDD5k+QSajUOG04cvRYwKY6fF/OK2RjTYpMxZtz7rLkFrSEuNY5v5l8H28QlxKp9RsCKuM0Oaes
afHVS5DWrDkHmt7kyRji25bJM4KyTu7w2TV+Hr3IlSZdhXs/DGRRiNC4JTLo5yBQde82Vh+NwxK9
+KaZ9Iog6Ku/hQJfy2ZlFVv5X3G86gZWxOJeJVojE0QpmEi3ZR8GhC9mQgt8G1C1KGbHSuw+9UsD
ltIs/0Gup2syxsGteM0AJ3hZzcZl2fSuFTsNTo+MD6Xw1XYFQ/BFgbwRi1I8CHOXyIN96Gdv+k+s
dkhHkB5Um0MCCBdCYt/0A4bXGB0W2RGWdm7gndZ2+XPq8PJ7iDhhjqooLCv2fZ019iBcaUfZgjP5
qtYHycUL6Nk/LXm5be5MG60A/FzTQ9sZQb1e0ndW5g1MmTVVXQTF1MtWSCq0lWaFjZwnrwaQOedM
ipfQKzuF9JR740DqJqwUVfhM+vah4/ZWfCFNsHMb/FNEzu2iA5T4GBAAoDfwt3dHKFHBhsx5HIvM
NP9xfQUWZskojVGXEvlGsI69H7p+Tw8D8dPIx9451lF7ZcHf9cUxAFe3HxdyowXZMo2SXFzUsPUu
FlehSLlhI+4aUklZSoJoBn9fHW1ArAxrVwutGBTn4MoPdwK0IbKIwiyXk0wW4lXv0lnzCS8/T6fs
WQgWOfKeiuIeQjJDAcgZXZAEhs1dbR4KmOZ4l3sy9HKbv3VkH6zatJDLRn0GxAjp3y+go7KDb6fp
uTiPwNqtDZyf4HeYNetkY+shYojwexeTuXiKPhzFEURE7bSNVJavD0DI0NrWx890WEv0ZVeXNUZv
qUpk6YT0E0VRYByyHpZPd+beYpeFD5Q6g0N0c7itVRknHUdI6VS8TR4M8Y9w5/BgFVg3qZXDkG8l
1gj+FkUjtOaq4fXJlpi+ACoXgS/YCpXEFatrGJUzgXz5cKhQcfx2gr9nyeC1ImWb07ss/UjxiV94
G5OKeiDcYNSXVc7KoyleL6lT5KvLBzxEPhrZO3cf0NochcXnCVAgY7piFVHaTlmOWGwub4xwWjHb
lEVBlbIQ1rRrTLo1rsnT+1dzKpAjocSW3rphJqkizPPOTUcjxQJ7h0nd7GzASQ9JRIWj32onWh/z
7J7fHCEiwLAqDdLhHkryrp11yryk1L1Y3WksIRArSTzkABjek9NU9EvfNa2RgN5jznWwQqkg15ke
8NmAx4iak9Vbp7PBTMgFH8Fc70G3z/9laPKI7AhjgyrCVhgh8Ax9+vWOxBT+nMgL4I1lH6L1VgyC
nvui9QGuYjiY4QT9iU5k52uvl/Erx1dxQSnKlNJCtYB/7LRt80NO49pMdKd3rDTBpkvqc4DvbOEf
sAzSOmEJ74fbclQhCn9bFGh81pzroGt9q30aVKrWJi+TRHnWy4SpSwXr49S2Vt/uvcFxDB5CXudD
L+Q3DSKPsP1ZkrQ4nNgqu/dKJqpDBk/8IR9yVQ4HAXura22+c6lr74XhjpBEazHFuAyJxEqTkuhu
AVakTwZKSrKAn4gSkRON0GSgxmsZoBG+mIIcYrAQVBSpyQbWfTlH+AY1pfck1CAsCyFBmuOz3Tin
8V1dI3x9Vx2dr94LniCPKX4BKCQZo0RRwPnIMX6df8ZVMNADFDr/wD8xMBWVM3bmzHMVGh3aFxOG
3SJAqlW6DIAoYrG96FFf3fV4KWtmno7KOC6JC7gJCVMd6mW9cKaRZrpbh/ZRFiNZJVAv9DZscRln
kWAWsTkYLTqS0w51/3rlfLXWweFIye2gc07qRd3gGSAlqNsjbucSLJhF31Le4HUztDqu0rJcySVv
iOyuOct7QjlVZp1Ug+jww4ivtJNfbDde+ODJbIU08LSjULXR/GAPmxM1qe3tWSZsu9VX0Jxt99Aa
PtjJD8xzSvvJwE+tIt0iW0hKLB9ts9B1oAoS5B1bhda9mnRZSs6PoTXeDB43PZ0dy1qr3sQe9ER7
DzMMpoloDKeyiJjKZf2RbxdEoaSk5wlYLG2TTEVlx0OOXTO2FtNJL+6sij0MVYuoVg+PJpHwzuC8
+cw812Ufi6rPsCceWbQmHnDC6LFiMXK/0scpgl+cvPIylzg5odfFje9W7GIHX87puMww/pQePmSS
SMtZMxwSUQqswAPfxDDi3ySPdwysWu8gUv1g9PmQ+Hk4RfXPMpZ61KGchGCOU6pmKs4JGcYQirfS
ix5mwpXFrzaIO6DDc7w18ajXyd2dYsw/qaAqtWPIMNLDEUrGx5rT17ryaOsyK+eJ0zVCBr0wPI52
VOSTbElSGHeAj0bATi8VNEtcKu5O4Ava0cYooZokgYmmPfFHMfZRwnHqvVRKbDTYZU3HhLCe8cYT
eH4QBLiRlthPFa3zrZ7Q44am7IDECiszKYZfqSjXE/+ZIBGR3ZC19EWk9IzEz2EHDGi8SNqKsz0o
kyl3AB+UmCH/F5G6nycXRYC3glrm7FOSJ36B0bGpDxUt60wdC+O20DnoaEfbQzmt4mlAjpwYuVVI
lRejkPQvDBV/9z0/kYxgk8HqEdRyWETb82JKjQtHEKAJ4vkltK7SIkDbo/cW28LY8HSrzYtdf0XJ
rX6F2cM73mD265C+FFfVFAtwmUckqmQXL9gLSzeU0lwY5QrGJ5ce77gwxB7VR3M4C+6UkMNHTncX
sXYYu/D8VsKRwFVlw7yCWs7Mqy17mzPLmswkCVutHJxOvFRVuFuNOck1d8P5xh+3xKnt3PZVQFDK
hkI7m8NvorGTn1YEUnhwfydXtUbsGeK382O7AjxO2yNARdV4jNMfvd25or5WyGt5ppFcb6TVz4YD
AvvNvcnlWiwOYNTa3QMygX3numWD8UzMyFs88PXpXuo/hfj2k91VyZi5U5TolcFD54MjkZ2Lw8yk
IzowSg5ZdEEA5WTSLODcPeqxpB5a/YnxoxBTlImQ/dCaWRlaoR09Qo3D0iCK3mwoyLT2vDqAZidS
Eib0J6Tv4jrbf2rVt1mrLpV21bU7SZTHvC1mS8pgVqykNxg+cHVdos+LOzuJJx8RdgD/OP3VBpB/
uwX4ZqYM41QWN1ohiCyAoY6rJ0k1uf8UZ5g1S1/MwEJOoOcWP56elEvCTZSWf7S5ZYoSPBL3h2PJ
Ti4IwPOB5g+gTy30ts8Kaa+j1HwzISi8X4bVbZUnIlWeVc9NliU2poME0cn3n0TDrSFhJnwcBt6w
fVCVJaf4EcpHbbrIsR1h7GwmRR0szNgH9iN9yLZsQvuhqVuAv3lmtrShz3OWCpiJuJNDIyfUBmq6
lapo65pX4pcdOhKrslZCkPE85n9s5TUnauLCE5O9BVyir8YpZn44JKGqQejjaBqZ3qfzYzwqN7Bc
Ku8d99FrbZV+YqqHe/eVWIXiyDTt7zqSV1M41XTMnXJI9bwPt5axq1o5RD0KjB0hcaTf1UIgXrVo
6x/XMjFjbfjXxy+d89PF7q8Q9QKfh4k1rtVgZEyzdf/rprs/cJS6Mcdam5YObOzXy1LUnDfcANxi
t9E4dO83xuU7Jpngm+Cv1LA+HYrLeC/yoy1sGBHYH/NtdfOnmO674ZNgwTDWLugpgtod03t7cC6b
w9ZPlLYhskPg8wsEzGLaOIJHnVk2iouwli2csLz3BiB8AhPLrpUO9YV9QqQRm9luqkRRJbxpzjUC
yPM0SHEOa+f8cE7zeN9jp4OqJSxua+WeYZ0uQ7veO7pVxm35rM52UIoKnp/WSXhwRw4uZU+ugTla
I5ABQEAkL1SaaeDYVoLBFC2569zDzayfHFcG77XcNxv3ig3eU90bViJXVtIDFI1v3jY6g8R3P8Ik
8fsjGLCzRyhXLvvwwXJkS1zRHjpJ4XQrcicsVv844oEy3NJ1vKTJv+Y23awHuSCwZMKtjIjGA1QU
wHf4BD2tXcXASicOdVA9SUr2XfKWdeGu0kFQiXS7prGM2+c7Q+vL2c1fDh+9yMNJJfvgM0E+lZFp
F7qPCtaDp/b3YvgBqoCteJnXJaPX9E5dtiuQzvKil+XAe0SUG3iYJt12Fu0JCUUDIqHSpYTuNKle
sMWmjClK/KqbySUsve6NVx5sAHoge/J3UNG8H34k1Mptu0i4f5NdAwb0KvwLOPHMKcgBY5yuQETN
GxrokqIOrNmM6HKG3DYyzjOckqFuXIbgXPXFVzytSNVPSOWa5+1B3ARpq0wGniVYxX8hA6AFMH07
dWvhzZl+B42wclRGmNsp6964+B9BSw1aGMekHFBLRq61YsnREwh8pwImh9bzpa+GPxZ675nhLmXy
SvDXhGleZl04hwiG+IwAB/lCE5KjysZ2aBYQhRmdxaENwdaxmjgW0TtxJr9HYJPQPeNEpdTPyvEm
7lSqbcBKZj8wYEb67W0D48i1u2P7UkHJ1/xPZvElSToXGLYf91Xtb+/pILejll50j522YA+jq45f
g+tjRa9TbR9wmyxTJRf+AIzKr9tPhYjFahHDHLAfFjOKtJqXvj5zvHtfQrF7Wf2JDu/kUhVgRQp4
tvM6SxPq/P8sefFfSvrOonEO+BunYHqOs2/x+FuQskcLnVKYHFZoFUADMYBVJy/mPDuc8X5BYpo9
pk06FTuAaJoH35IKg9kDe80xM3lBbV5en07ZH4Ylv/+y8YXe8TgPx+n6xvrGAyG+H9A07dbFoDjO
DnNcEkLMjrszKna0PEhRDz6hIdfNt7baw2YCvOfzs8RLl6f5cCNa8xaWsqi4U3njSS8TuzRAPT5j
2SmKG9Ru+7Bv0MJNRsfuofoWVO90vkzT7+yG4KvYV74X/uzsYD4bgv2GB9XlPkCNshQnxWMeD9D8
TZ6K9r2dwvUREjDKLATdIu+S+6R8c/wDBQnDuCwwhn2Uk65S7073Lb3/iBrySgsBuqncWbZLL/qj
+CEB5SGPCeNfIW72jfd96VGkVy7aXDNviTuPIQe+Baz7z8XbTd2faUZJ0BJkkgtzfcY6Y8Atdmty
D9Asg8ZlDXtJinm8Qtd6AI4S7HgF4omKxmBMGNZO+8sHtOHL0t4+gGR/5Bqr/gJNUsvtwcRhQn4b
gFN84Xt531fSSMj962pZZbWkR+QG9OtTb1FGOXKAhuw9wFDrKPtrjcLDKAij4BNZ/ccL66zYVsFH
ItooVvnm7jY24iEVizdlHYZLVy73mslOWmMtQNiDVzk0fiOYCxNkdgkcYsPQ3R4/7p9/yWlDBWAQ
qPJo8QY7iDwZrIk6hiitH2y79S/BESmXu7Ri/gZ/yeQNNjJAcE9cGK8lQiIjNvs0l5zvtFL5VWE9
olePaIDS0k4F6JW95iQvR9iYMb9zI6PEgVzY1EBbRRzzk2coL37PPNPO0OL8dAu4PtqGOQcj9bPl
kJJ+IBXWQL7KnMYh/rujYhQte+1jFkWW+6q91IxceOfWdme/nOJjBC7+OGGRaJGrqjkjcxdgfJaX
7bt8wm3YCl+7/E3xsWHx7cfWBlesBr5dunNBRcl8YkzyMPlP8RazRhASRxp/k2Goo1G2SgzK7K/4
ARFgmIUGgQx8kYn8+7mz92HcGNWORGQ5hslmlJ+BpgRcdOT6G7TPqfc26SG8gD32L/mioVg20nT9
SeWM/f/pyOl2gSpmykpepvPc6Y+XP+c5CTnqUDU7JKKG7iCbhtzleI4S0t9cmd6UoV8gKggy3HDO
K8ehbH8gNqgoyMBr+DcvfahOODP9NATnBZlAVGKo9mUJ8o5AVM7P/8eGtjWCxkLR2s+SfDzXIs+Y
64I6C1RaCxWxseNkjvJq2zvmby0y87MbjDiP8cWBLq6rPBwua9ColqJoqimppjQrks2VCJC/Q8ih
6K9UZCgbRYgYGy5l0mCR6kINwfJgjN8PAw/dBNnUwD4mJ7QM1wM1KWooqZwLVjYvm9Dd2g0W3R00
z3VdOvSFyElnAxXpHpKOnjjLYEpIh6gkz5kKrQp3dzR7vcfGQU3OFJkvc1Audisp4gVSzmvz0PaZ
rAbPSA5TxnGXEgNEgUe5tj6OrcNThV5RhUgWSGE+HBzzAvgs4f2dsmrzWchDjZxw9cfDpbQOJeKf
Z59vfYeP4cuFL+z+11MFNNqu3nXqLqAfUAKfILzwiLbu9nYCip862AOumvY7Ymrdh5lQB30FoCNF
qi4QH4rgsW2SXmFcUK3TjfhrOAJ1iSf8cXGK2OyBqoaOyCOnGXxQzPvMFtHv4qQFcQZz4/+7Djay
6pMbgaCYjnSZn1KpUBGkkOSrYvjmYEftw1x3VEHMGpgwFPldJdZ7Zlbtsb3xtmeoC1Kc/ZUImKXO
GCV++8bLhiXwbHuHjxThNVQ1HVH7to0l3dxoOGBVhxeeiXLRikIqy48lNs2R/bmoWmsmMXTPP/vK
LSTpqNm9LEC5Sxhmifh3q7MB6E3MDHreW4r8bxE2I53Z9hK2sk6cBXqA88HrC/7Iw8WSi4qe2dKu
DbsvrpEOWD94bq2mWrlYkyKAoTB0DXn1CsynrNQKyK4b/w/VwX/ADjyFNlc8vAuj9HwWSjLuyigC
me4Ogk76R8Z86+mL6K3PM4HMjgj8+L8GFsVN1p7J9ZoW+pPdFvEM1dkGHQTGNs1FcH10aiyY1pnM
9PIXVIyECXVduX9t/VHpsGjtWWp6whL3AQ+Kg6eGK2FQwgJZFU833IXuNmpBSaZFGqm2fYUCdmG3
euHvwrknPV4xg612Bw+Z/ePXq0JPdlhKN/nZVm3SpccZ0gCS7NW/peLMSN3aIxetlSlXsOeWuu4U
ttfWSn1BAyBh0uJihwkNarb5iOtvugEHgf+2DcGNL8+SDsNhLTP691saflwF8uOSu6vGu+yKMnzO
ZfgcW/O+3rKkIhfcgnTFBjsv3Iaiwmkm4qt8VkN23AmCsdtnu+tx44QGmpSLDa64msONzC5U7YVs
oeq7PvjZdaFDJpEMKMSjxgmpPFPl0qYVuAanlvuBGfNJxr9zBAdoU7GBsC7BShgIYQcVxIa19aIq
GUdOwFfUNN3xtuH7Uf4XizEHLNOO5L72x7FNTSebfdt1LOEo4kul+sD1cCUXS1knSR/7kK8NgF+k
1rNKMV/l1lazvQZwR/nqsxspNY9/egWoe3CirqvRrGMQRE0ZFHXDjfHsq5Bv/xFL2ic5zqwIz+Uz
80o7K44BZBeLiyRhjdpwIe78KLay4ok92vd/JgIjDLQae0z/QMoq4yxQtSWJgUbSqlabmsuQcucn
h8FlS1Dj2mYwH3tunLIhJifZe/91opptRfFswQZJwS6GpZsyhofWNJe31XYdSV1QKiracXkR+c63
K9xQY9KhpSsOIpZRTY0loEVCL8OuTQFI0Wv5IWL0cPH6FIFZYYZhWhSLveTAWJmp784bw3FzNw8t
Qhd0bNhX4Y7jx15l6J2T/st0gvOlKOPvbq116t4+beu88NGZqsBvxsSnagmvdD7HbebRDa2hSasi
ZAXvV3nYK51jGiyiAdT9Mhw34p7jUJUKQPIGlyNG9Fcmerw1E8HuUVmdtYEofWEa4t7quW1BHGLr
x6VqlerehamtL87xcRGZwT9KcLjEkPoSSBatKvdxt/pQE3qWxb/2DYD7G69vXrDn1Wg/YCTXtM5x
NP+3ubX0IoSVsyCs5HoWPNr5P0x7yhzr3qCNQW/D3qNZtn0/aqm7L6xSHGw7Ie/SKVWMlt7OXynf
LvgTWmpKHOKiHXuUyKMghTQNbBud5u9rQZWdeWvcf4ujycVgLM1EaZzxelN1oWXVHR/qtnc8clmN
KPBwcfEw8Tou/YPPbC91rk/GJSFo8v/ouebzbS0dVWn4QjCS0LKxb3kUD5g8QGr3ghNlJ5gTbFVm
FBWfezCEiuHrtePHPD9xSSXy3CHaGSpAjq7j6MH+/gspUWsOGFtODnrBEkNt2qEejX1mOe9jsZ3F
qYvuvIaw6R1uvaL7SsVXfJ8by0hIqtBzG/h3lk9zL8c+U0F90Fr2/ah+oFw8lLHCWSLEvUKUFk/r
GBT2TMWMI5cqm4PH9HaoXZTDd4f7PGs9ssQGT7kiOTQ8nvnMeAl+rkooz3DpCls6KdywTyNK3WpQ
64F8pXfJdORdy9NJCI0zCIzcFgoEq6jemgb5rwl677DpkYuGtQLRKzmRKuLPYkp/AEohJ85/9lnp
DECJVLrSC61WqwTEUQGcMHzyxZTomCicFQCbdPQeGTczLljCsaL6JJA88oYINm+1cGEgcENir34F
ky4Hg6VrXzwUh+6WlplVXMmaRkkUJIi7180ex1+HzONcIpoFuiQyw+zrOXHEwHQEkRPYCC5UsHiS
CUT1768B8TmymB8pjBZsI1VQN8cmjT+jRL61r4a7f1+yaUied49sU9ZGD/ljHlyyuvhcTzPzp3kT
1E1xdz0l7dr5P0DMR+uYmMM9pRgjznJ/qnPFuYh9PRRTQs826efQRnjZmh6BzjjSvopxBhxp7jqh
d3v4QX20MTTX2FbX9CcqeTsXoUtFfyy9L01ppJohEF75bQ2HO+j8gk5ynmd0uEyiCPE87JUwSUSX
PtKZORnvxVE8UcyaOai2WXwnXVhvG3TnsXT5UKI4ddqBYnDPisBlN07s+O+585FrA2dT6ypsYXc4
Cf6zYDWhlZG6qqFu8DWVdsQlXRjkmRcW29vwTeQw27PumOZ8nOjnKP1rjOE0MxxP/yhZZts/Oyqz
CAYHL4+vLG5JFvbzJ6eA08BZ5aqfteoCRV1mv84zWnBwYe3Tbsbqrum1LTeya6KHLALMBnIAphf/
aSRDd5uIW8QURMOaSTLZYtY7GA7/4qLrsfibrEz3/YznNSMjXLRCX0GlJ7xOkGAmMw0FgJj9uy7N
8yqE/l0pIHGbhTootvJMRmakqodoF4Fxx0PCYZMHQ/lahbsFByNpxo0ZQULA47Mn3h8emiN95HB6
UixOTQJ66dRfaKgMhmZYOHEeZrGm7vea1A1rZJKWU39pgc+IT22fphLMHDFOrbMqJBtLZg2qfhi7
Zr6SZAgG3f1aZw0gtHYhY1cZO07GfGb0bRzTfpQTy8bmUp+sBItlTtJOFaCZVcs3D7rVT3AH7711
aG5tBuacNMFWksoE8SonUmd2ATqB8DgvC3wLm4b18mZjWeErjGjP5/VRTG70tvMskns6+tTirnz0
H5GvpzacXuBqHACi2i+x9b9MRD71IuGFdAUM5q+Qx9F38OgaOVo2O3PqsxX401cu+VnGBU/H0Plk
x26DbEV2Fv2gthn2eaG0KC9426WF7ifRmyZqwmQ9lcaHL8oZZaZDobCR5PlSbnnnRH+WX7i/rsw0
b+Bx4tlpk3PWR8ukzF87XT1BUBOxI6Qt8Byr4aatVdG2kgSerbf0Q/C3iQN+TPqfGJqoTBhrBc2c
HZVCMWbIYT5XZM2SBXjV10ZDBrz/lkkErpdL2A3GGtBZuCtG/vsYBBTYwO8jMZwZYDWA6H3L3+bN
3WD/sgOg+zkPhyNeoltDesGP2ISjfr04z2bBRBlE4Fu5MtL4ATM1jMOk6tBUct2MXI3rjeVAcaIe
DcWPXNwgrG9mOGJI/R8iykmGVQ7Jt5sD8CzzX3+3HIQcjHYTOwmXqLs9yIqbLIUp/f8tAApSTFEk
oa/AEpHwoDUpxgEeMSV6fF0QKZ1zXMkegDw0W7kbSAHS9Jd4ELAn5z6g9mAlt5jHg75q3kOeZn0B
KUmYesCqfkUyDmvOe1HQKZPbSZUlLR4nTLed7yCVHxdrfh2yRSSrjK+A+FNb1GB4PpJ9QGPrJqP5
VhYyLWt4Nlzwvv1iVErPwlNbIzrrEA12tSiikgjQTnFJBC25KbGPUm36f5FPJnzkfQEWI1QnAUOe
e1IGvpkE8C8luVWOPuBWI5vAd8wWsfQmrrZUxw5ai51eWdXc6kmR8C0IJCybWbtGJQs1ZAtPmJMj
vzSbpMsNO00HpOiwx0uIav15dag3RLWCvkEDiGel0EfdmP4p/hBN9DQmOwDktwBWV+eThPxMVjRy
i+ryfffrMfi+y/QhJ74/RXBt25pJmBpr7UN1cwpYa+fdBuR22knc8RrWnCqELX2BQbaVWYOr15F9
HbssFngRJcn7kPeqn6Xe/kSWnyC8/cd+/uzKCYGKRNzY2pnX5paEcwVrnPVlo0bNmxgZKZM/hbu5
6fgQmoiPVtmwvshcK6HnhB29pnqpAGW59ncQ6rD6r1TSdW4ShPr80TWj4vxrDThZXI2Eeo2LsAyc
QIGS9boCU+cuXh35nprRryNJB0x6sd4K6G4jPKaTStBnm95vZ1641mY29ize58U4zQ47RjEbq6uZ
T1NeGack53SqsxB70ZfhfP/04CXU2LgzGKe8bNs+5jwTURuffaMkkcbKemqOhZJCt7bbEPI9UY8m
Fd9VWW1dV6kTuZ+UlBn4ktG91YHInqEyqqra45AmlzpDVVYhxVp9hWtlPNVGNEyTv/7hg2pdUC1x
dP0dvSaVy6+Yda+gkyC6gDqDZirdhO1IVdoDaKd8bpMISReW5m/7KT862KmpTEXmWLMZh6rXL0mh
9sUYGlXDdBOVvdAgiPbabFRPoVaeBvtYpSIMiyTRVDLBNn4z0a3/mcGO9xxG25q+Cuy/jUn0Sw9c
oGHopq4RJfc3lCLVvG355XB6PkTSSSHhmSPbrCbdQ+Xy7rvf2/lCAmxdZkPb69bHUbMeTOQJMBAi
4addAs8wAw6Watg9IZejKKmOG90rYGm1Ry5K7qA8iuqGUh9UZsqL9JIPOYBE6LzTjZtM6nVSNnKg
+wHOk/BlYjqKPHAaajavhCqcQcZQtNUJTJwhVHAng22gxbyngw/dztDiQ5MUC9jb2X6tOcgF8O4x
HPc5xH07YJa1Yfnen34plvU9C+8tjgj8KF8Gzh375UsrjIW3chtKJBrjwKiX9un/UrFzdn8bbuu/
iobHA/cqbdgzEfbfOdLA3QEu5lgLwBWB78VBdT6vIdfl14PgAePot8mcpwDJhmGUcBYK4+z3qzHv
DRXYSEzK+h/63I4XCLcmSANn1TzOPCX4PQKCnPO8iT24ganWSMm0XLsX83FCMibWQATEZ42POqh/
12wTqvEgtl2Uh/ohJaA7bUJovBZs4TexewT8QKF4O/ly6zI7iL9ONN/Ll+xCZtKT9RcVTCVPaUOV
rB7vSEa6/nBcAB6MHWkoQ99Ym1Pvn6Qr+E5qsxZr8zmauAKTBXAkN2LqqVfkQNHVL4PtleWZgfIJ
dSqpgUNDgn9zBHyBS8DES3oYzH+eRbBf5AkUsC38KLnz58hArC/iTyZCBBno+Zbn1UJrQZruSlna
Yn3fFbLDTBYpsDi5iMTLvBeC19sMBdENUv96IPx0jSDxTBy2+Ah85QobGOF6IOrA+eoDGVCopk+N
1utzXVyt2yFe1EgNTcK1Wd3YuhEa0kYcWeBrTXCUMFQfUezuRaBI6FLCq1y4SsT4F6zrAmyOTLdZ
SY/VbEIcmvoZXUXk3IHkCOje8NsDaD0z/Hqm3jSUiMn8kYVotxN3PhB2OMSg0eNjHnjdTsLFuywx
dGyGu4ZxSeghLhNHS98hcWxfqZGmbqdw+x1uKLmRpg0HpZuKv0qUWBjhfzJb/3ghhmCHNrknyaVf
mqAG+1GimKvxXN8Wf377uLXeKH0kkN6p5/kGx8x8XpAugsgp/3Cwe4yiZyXkq8kzNSkPedoH874R
jtn9SJdovf9Ec7E6cPTq01/TQ8mF7bpH3ViBH0/2Ab+fmF7FwT5yBKWPJArDC7kb9wF5vmaOXtbC
FJ+azsQl2YkVUqCZYe2RXOYTIikEkRGwSxUcmN96IZVuvg/EXU9rEJ5zhFBQUNaYAWsLa03s+i4b
NWtG+nDoKZ3YFT3u27HOJqBeKUuA9upfaFgMsQDuWckBVXIUlBmmVYlkuYk11RJXNUvQdsLf31W5
4/3smtmAfxESoZliov9FI/qBozl/mxHyAimFKNHjJqeUypspLM4W9CRjxOUCzS4pboFk8yMXMemN
wksiVU1uIMiVC+nWxGOBNW0VHhhz9os08idJl1F+k/AC+JU+qp6Ob9TEJLGjTFvXPMRzO+u11mgn
QCTubPvR/hRLYtR/jNY+IdBLzfAfe6N8gUyhoH0UifFekkpwaLsK/M/CO+DpreSgqwJdG6RAjLcW
3qCnZ6YHDZ47PrAx0TylkM580op6ZifGJi66MMUrtirx7rnHSv9epMaNoD7f27m7udzOdgDCeEOM
Qz7l5Zt3vPo3/FI/2IwKAMwU1aBazESfh7bltH/lac87g/R0F3+CsqNP5FTC82nX4L07rZGFw1zN
vtCSxv53Kjvb+TTBt6DLp9GhvgVt0edLzj9DYrI785K6pSHr3in1EX7OpLr8rB64R5ovuXwaV8Jh
/j/BkKAJIJHOMRrNPibYdcSPCXcbmLMiKYssS1D9YW892I5EaTWYZOa+vOEcnkw9dp3l0GYzBg3o
+rEg2LzPvDNhY2bJW5/9GwEYO1U/CaXuW7a9m98iJZD79zXJ3oko2gVJjXWHT8SIyOApNzQ3PzFZ
pNCv0YzZ3DV5ZqJKkNzz4LyeHiWXFx2uFuwt+awSv3Q+EJDbzs7+kkRrV0DiSUYQ6T3UUE4AjHAH
lt69YW/lrPdBPXePoTnAcRiheAY477VERN5jZo2aX07H4m8CN1qg6CsSXRXjMWAsYwS8DA3UUT7X
zqvFtq/546tI33XP3rqNH7cQUyV4fzxskql5amn8eFHT6BmP83twRtznfDLSRpAsNhmKdS3OcvtW
S/WSUUxnT4cQWt+z1DJBTtjGtsXhyRxE257QkA/O5PUhPd5QV1bad7KpHKXP8tAIVw6HnAoula8M
adVMmFWM/b2qmCVX10QMALsSSyL7G+wNz7OsUO3/R5K9HPurWAfvViFjyOAyaWKXz4lcy2RxwSkb
suI4qretApjhfTXWjYat4MDHe+lY598S5Qb614AkbgxMQd5fCwwyGlaJzOV9PDR3az2XmdNvtH2i
AcPqd5dVfaUCrGIHAhprmhd9Y2tcQ5IqFsXTICrBkjXrArdb9GKuk+Cq7F4Ag9AuOAMepKdDpDay
MTc+sAT++Ik3BCQukj2jRSu73WLBzQRoXLVk3s+aJ6NqmJkH7WehLFnU92Abw0jRG+XwMytDyRwH
gaukAf9V8NM7TTEfhuKUT9m4oCwj6UJ6SZbs+XXs4ZH91fzHWU6fp8ccbo9yG0X46z5UuOAh10vR
2/cfJ72TLLsNkpfZ9cfR8xC+yoHGk3p06RLQYFYmxMGmQn4PsxzI/87vK912gRa+kx1gIzGpCKau
L+MxuLKsE5KCapclzosmQ5GUGOZ/KpJC1yvGZt3PJh3sm7dCfNUNO0HGnSWcEpPdpE1Dp/NIVH+6
YLl6QLtBGj0EoPvG1FDJ++s2tFL1tWCXHM5TcF10mlWJJOO8h9+iv9iyPV8Kcx3YXIW64BpkfoNl
3YltDtDGIjM3UvmvY86I+x9TBUvB6utdV2LZqLIvB4Y3x/OdXH521gx0mQhKb2V4Uv6u6nRe4IJE
scRWudTpFFJkS5yVqBP5FzzkzTPqQF7M7jeUVVy1kxugbA8cOs+mbtGIXNzPV+YueXRGTzvxOwd2
pkg6r0K3slkvTMXp419+CcrCWHIJLQHRUItj5gHRGwC9uiWmMy1PE7psdw4tfsP1+FxmJDkXFYxa
9KuYt2CJB+cj/SfiLgcwY3qYMvKWiupC9qWjagGMDx+x1iJnea+C/i4mi9M2i3qcBMITFlcCpE32
zbNoK8hJsF1yxmRrU7VhL6CMnR9OChNigqHpnjMVbM+9mYX1Cy4WQPtiSRdVSrURQtEgm+x0pmcf
TduP43ZR8wSEKke6TBGpGhk7uonVVcwCavObExm6bvofdjZF8pqokxBAOTWuNAemyh41DIX6RIst
rL3aWuII6UYj4XRVNMX3UwTWX7reiQl7Lp50XswEJTmvr5i+r0XWNXKTnKNhT03cEt1qgclvfcAU
zHOwSAPXGAtpOq/4wTRCIJ+VQvsg2biX9htROHyOP6ffIsJfXsWgZgMOl996ugNN8Lo3wZWT4pvr
HxjdHZEHBTXjdm7bNc//j3NboiGtggl6fU7fQP7ofCn6pZ4ViDYbR9rBDdgxCdKT1MFXW3xf0n06
dYwDgs89O9RjzdDeseoCaU+lssUi6ZPgWkD0CKlBLZnp7k2ewioMWrJQJjrAWBOBfw/DVqzEUHOM
2ZcfX1JDZFWEvb7365sfFnT1McdWouO+z2kBKk1dEIxUA5iJWsTpQfErLt4A830gjjgkT1CrM7gM
DicGgUbKaxh+hscs8b1QiaygTI4+QLzGHXf/QL98FsB3TPIc0QDLpj5wh+EBeO1b8/ur8rz+fDKH
WTotuvw+soT3EFjzfTloDCUdRF/Z3baP/vODc9b/lMMky3t9H3FmBuzaIZswuUFq7pL7EI5kcNPG
/WksYmYC5WOsFbcw9+O1nXgMUNB6nMO2HfBRXdZUx+9RC5aKVdpj9mJwroLND+gDOOgweOkVJMz2
nJDFFuCmBX1jD+wxVr9KcdI6V3Zdze9Z+VKJF+O15jgM0fFbXcBBT3JMG3peoDN5odJe33BKRvXe
XmzAlyzX04NG5Fzl4AiTxrWaGhfBDa2Q0z55FSwonpPF/NvuH6bXfntU98NoknjPRFsrslRbcFRg
dkpODf9zQy7Q+fhBiUYoECM+yFUcZ3LQb6QjAD7TRNjKcZNRPfLMbxDJE71xZDJzZNmRbYwsa7A/
IDaL3hRZCZGaBBRGZ+3urbREHH6Vo9OtOx1crwP4MzVYWMO7+6C+HBmazdNUTu+E54tfDqD8RID7
M7ZAhTeYqnkZw4ThwX2aHrqFbdbN97G4gm3x7iLKwnZStrcO4xocC0dbaAOxG/fxI2d+UmifrDgj
fM2GuVGbUBeKXiG3I5aj4AZrzZ9BzPhr/UGm9HIeZhvZTs3DOJHeTDx5QJxNHgc+rPN+n7uCZjqJ
ahnjOCgGWVsJ7Zzh6hU9HyBkoB8ys70XdI+6D55jE8fx97QXY2QAP/jxtIEMDqF7JlyDZPCA7kFz
/xY8sq1WJRkK+G4UjsQ84MquQbmY+C9Rxn8HbcpQXyFzlY+l/bRxjq8ffgUufZw6+d46haOIKE/l
yRIZJHhzixtoSfgmFO/EmmPwg6klcQxXrCf86tfZq9bMzNXjKEPJgRgVNCcmyO/iixR32+m2ZFsO
X+/d2JzLTzgnmxpdRXF5HIwLRZbUhDYkfNxI6+ivFG6PJ861FFVK54AHeycjcjcQOrQ3PpCfqZOe
/tZ7KeLlAH+TxXnWcwYAe7o+tqbHOk5dVrniNfrDKFTsAFHPYfYrM+h8lrB3MMWAfyKY2MmSMgyI
DUCDuxxa/hwSuZ1hlJh4mkoV3Dao2LzAhm1gGJqc5mZMHpZV/SkQHR+9ccSlseUb5ehEGU7epOCK
EhmpAl/L8cWIUobsA39ZTUGLGFpKwtOwE4ezAjHMhdGmqCG/QvyIajCQBEre2JFKDlkJ6OHxDdPk
P5gHsBhJj1JkpWRiUcpmAA5nUqqQ0l2u0iwQSVprY0KePptDbWU2md+1CAXYargs/DhNWCTs9l4g
uoSTpZ9F3e0sq/DM9XvkynGKrReh6soaS9p7CDy1zF4ylAc7QRXovjefR9OrgoZXGoQswCRBUQhB
Bz9untQ1XxBnbd1Eo9mmVwfiXa3nll47QIUBWN1Wxx705jecUKfbC8D1rGsMW5qTKvSUdYJxSNNf
/OUObrmJ3ScTii+qpKT3K5GP4xmhM1Su7Mvl/R0DeHKKF3ujNRAmcrny+oTDYfjBM+g8HdVbvQNL
emJteBOqO28jz2YjuWDz++nlFO1ciklEl4MZEa4RKRKkKB5U9Wq/7+/WobxkCtT7baXSa4dXB6RZ
QmrSUOEUUbrlz8M0CiYkICj8mgUtAGfZkq2olWtIXfefWV60XVI6tSvulKIhPNw/D9dmMXv4ZjCy
5g4S/hDVtMZMS975aSa+bDXSjpYtiFAHiuRI30+D4K2JpjWEhlrvrnUlxu+7QFV4abWK/My/koKD
LSl9t8RHluK4HQN8R3WPnChwjebhI2Yg1bXPBvwSR+cF7vDjmaeJm6bdSOjF2vWRTUbTQQO3ctkv
lx3CV/5ojCoJbjQ68k4Pr2LLepxKYjFOXkmnNhlgTGGO7tp2BHZMcvobndIDSkjSuAl2RBKMApaK
3sOR0YDuDATKMzwauuIg50M5jMG1lRGBI/9OFYI2Kdx/VsjrLzibUUgmaXjXTzivRXpRulDTQ2ea
DogXAbLO4ag5CcJQ61V9MFQHLMrNhhH2LhGEwcbIlPmi//vTqu6S8PgMONQ7S/7fKiOqvaWMkmKe
s6FQ98MtPyYI3m01g/89ZYrNj5dwnaIPJkOsh5/v0kbIWbAT1dP34SU/0i93Z6cBoRjiStmV5BeD
1/XkvA/BjhmxR+gPtMVKP4ROifRLdtfaF+63OGuMH8T+smPOyflz6vEUSjbPVDfFU0VyoRrp4xq/
JfLjVA9fmOvSSbkvSqKXp6S7vUgh/YpPguAfNK6Wwe08qMyf5A2NAD92DbPzIhZBt9CP+EK8/uPt
r1w9ij8Y8HdA0z8i486SuDZ+vQJ34ibqBEXOPhHKc7tCjnz30Or09uvHG/dxGkBROfx/bZr6cAH/
781Ja+tlhy/OhQavds3OnIQrIfboMuMH3pvySDs5qmQMKRqrNomtCVzOLQhWmF0Dt5vWcfKyVsXZ
GMKINlNPvj1q36JQass4cQKpA2L4Z3bbOIvc/XNC+VGGa3/eMj1FGZJ5Aap/xKSo6O69FLfgPidZ
lxLxum7KhUm+X/akv6OvRPJ6BAR9Ckhdaok8ERFiHgrMnWcS4kzkTZOVU917UTaXxFepvCz6ahPG
68cSJUgDa/DbkAHd0h41iHwOx1ulb7WxHJgKLoKxD8uIPSGeH+AC1m8fofqrRRMbPncrjxn/E149
d90nw988r+wNAgmoBQuflMpzRRepW7u7tgPWgboZwj8489SjJJfnbSZcn6ZYIp3Oxz/rL8i4+XKI
hZGjliADHAIUEFmmFMvbLwprNB9gSzBPknOcwpUp5xJc7o2Bj2UPzelNjhwQHEtjzRoXZTVC3LfM
xTxFR9cdXmLf1AX1S3r6hl8lqV8VWXqyp6rOimtLHs2FelT7LhKaqTQXSYUHX2smJu0XwAuVDZZ9
NllcSEJ7raPW1pxWR9YZaGSXMLUq65e1gmWi1+voFjg48JdE2a5hbTJze50FdpyDrTXza/pRO3lK
SG5lIKgfZNxbOau8omKhsIJLQFMYrbnSRgHTPesGRXJSrDkyaw9GHNucqaZpQU1wi3VBnkwVE4Kb
ma9AHbnkKoeVo9A2MpjiA/s54qzqROs50tYQn/2ta9hv5lx8MXN9E5MrH5DgxDGLLb4kXx3NzrgO
TZqlPq/bp4nYMToGtgskod+9+NhSKDiAuwFDwPQX/eZ/7RZ1uPkaI/1r6IhdyZ47k9rPp3lNc4Kj
PySBhe6T5rPt0eKZQofGn814QSV+8phmpN0tzCa/IR17agvJNkYv1L/FpBYO/CcP0uyTBrQ3Bn9A
co9l+TQb1R6YCpxhJnDQLcfp0hbg3PVdILKiOv41LJiWrcW+N5ubuTmaaX4+9/B8YhSOMeufGvrs
QBtBEq/jPQ3HwwQsnwSk2oOFMBO07O0RqDGPIG7uEDKN77SV/V/FgnQxe8EnQTAuBgm94yIQ54xp
jsL6rBYtLpIjdYqbN+3/f1oY0pYonKPtMP2OIdQmTTkSdQBCjgSwaumQo9B201//oSlHeH4m2ROO
cf7IhIYCmhsqJvOAK5etWJTLwcXdojbKy9Igeq73Cdanq2XfF0Unj5G/IMTu93qEwcz/PpqBsCj5
i5X4DFHKOAi6y5ycoRP10o4L9MumKh3xWWCvltY23I+XwAyq38kvFzgG2a/FqlnKbwLhOhDeWfDt
9+Qz5rukCyQuIiSHeTEoxNTXJofRL2Rh54rxvhpR07PZBKNWl5k1pXD+T1s94Eo3xTeh4EThdWQg
+JjDK7ShqeQvOZuOI5760R4P28GDJr2/d7Hcv7tHJxZT7exHgs7GSz+pEvyNe+TGxOIfLqoHEe5L
3LPDCSHta/7u+V180GLaQhOy9TaLtauRoVI6alJQoP75FYitVLrblqQc8efESqoFkQynt0e7DGue
ifBVVLpJxniO9MXxx07zHHtFhnYnOl2OiihoDBWXRQe53ziFUWdeqcIzoYo5h8d0aQzdpsQfaBip
8zVvyaW5Nho3iG5qTesoB4/R4JPn0p572I/Tt/7nDOiU11UlE3DHMBAgsmz+aCPJgYhQbCQpE/dp
qkQF/lAK+4gWSoitihzUCT9LpLIBm2JC9D/BIA5Tragh2/Ip8fLeM6rWf3laFijCW4SppwgY2wmW
+YvY7w7cWbVMI0fdsF8pWLPQvQ/h9JS50Maolvc7QnXWoHwE57MWf8jnTJw8PI7xyFHfThVZMriT
+IMWVN9l6HMaATlovoMw+OvyI/BNgu3pEMGqL0udwrE0P5Klc1TwGd+/aNeJJ7eJpozf2E86u8QD
qnh8IMe6JSwTQ73PClCKJ0iJar5PEmu/8p3fKikeuGM7xTUerdVoS5Xs9U32jz1JaKWs7H1CCYCN
QE2SFeKTh9fACSnMBmSmcaHP8mti3Kca3z2UUpXFu3GEL82skPfGuNdrBd9OSbGJ4arkfJURhCck
+4B8afi/9aObv4LpmFrozTdHLkjUgWr/1NJ9Zybt4xUWONk//nQ4xtVaQR4+s9QoX3yh4KgUa4OH
TBTmDj/axQ1boWSYP2JJJNirB4huMbbuIpkG5cdiqVYZu0T606L6sKBF4eiuTtFh++mpr63gywkW
onUpeeuNwcr7zyQWUgN8hSBkIznC7/oFPd3jVO6rpW0+YdjnzBEEwu/rGpOrZSBbIFEsWaWoRaRA
VUozELYohB+HO7HnZURVVx6+YnXB2+cQLSPnVPusLb2PZbHknCugHqgTjPATtsNhrKAQt/H8YB+p
uuOmHfQMiD+UOIV9sW5xmYfcdn2Ae2sEvsDn86DR1N9HkuK1otprClujAKAwSgcKotapDinY4kzc
LI9nPhYcZiy+zxWdKwVVaTlbHu5QGLAGJE6MNwESMFs3ERNCY/gNRtmPCYjovpQ5npUuUpzD7d3o
Qerhg1JLO9kN+4UfRymQ09BW4aPhlWLDytOB7RMmhGD1kXJGOICLbS6WwqTKGAVRV+JxvxOM8PgU
5X9xs/sfb9CjvcwrTxZ5lV2H+dRbiivutDX9Av4x/MJZdFhS0IEL1No+23M/KknPBakGtjoJrqnq
1yyI3d55f0buiHJgXt4K5WY/mNxLNy6YiwjGLSBV+mHDNcl6TM/7xMHC9XAhPEboklV09/Ik5hQV
gWiosfu1piqyYs55o4IZ7s57/b/tb6NijQ9Msr74PhFtkSRt3Y3KiUR4a1FDF6XjrVftEnhXwu2I
4123d4LwsVHRb7nz/NqS2u+FpZvJKDu5fRtAhqG7FEvFXqc8iTrBSUjMW/y8x80nA8WReCSUx9sx
X2lNG99Qyj3DOBCCpZEOvVA4BeTbOhlhy65ZPrzX6WKerkjbATlfKJauIlGGqAJre3/dZS2yukkL
LQM/YGynPcjqepsT6XwLIjl73EU4HSveEINPdd1z0E9XQUhqzf9utdFdM2uvwG9V8scdNCkfnfik
3BZxpaXoLGLy7j326+pEoVXtsebkHnhlGjbXsNA76dKziuAAFTVu5CBJfx3trCegsusESNJur8so
vojSy/wg1DHLR1X1kdZF6EZAJUST4YmAlkss6cmXp5A4UDiq8Fh5f5WDvx3vljp5VGXlMH2E2Qu8
jY373SFjap1HcdlCNOlwfWh2xX4ZOPQSU69c7aZCzvbt+biFDZPHGVRtvzDWGDSk98dGmwTPk0Q3
XjORd1DzNj+AHnMYst6c/qIkHIf3tjAdZr5ztVcLG8blDEPJWdv0ITapGXQTOMEIqz/LpBfdZS9B
rqOI/52zhcmS449hIoTllRiBLV59ipEKQB5FV8LWjxAx08qgpVxOJL3lGY2G7rI7M7ttg42NueKY
8PYynIiO5BHUCyEYnJyKzQUpvTflSu7OsvvQ5c6Ejl3BoSr6LMiuTGh6FwfVujvkuYQPzEZu814Q
iMgCRCwgUp+pSafQCkAOzc6KZ1oPGZx2rIAuP8Los3fwSyQ1sTcVWwlddaGFZnEPxprF1EQIVo7r
18zqwG9tC7HGzjiSzQMB9jqoyKL7/KSFO2M/Sr+qM2Bf65uHT/PHo2hcpV5gMt0QQ7/H+zPhOBtE
5b/CFa6A1I5atu5UPmDfde47fWM5q3yhLpmrCrJ4jV3iKbmPbERFxtKgbOCjROzv6LxeVpyRiX+f
9YqpKqb6xQL5HBgpOlaK9YxsS49L3IoBY0LzjzyrWgTaE+5HYhK4jgX5Cd8VElRDMPnXk+1lMkM/
i9jmB5K3ZMqhr/TuYzttpdpvAF2GbDxg4Exsn2kVjTwe5mjfYMOo+lDhGgXhUCEMq6cnVvIs65V9
U95sCsb+6d+rkp/jq/FENa9dekTq5Fp06xgoxJd+aoDT8jjiUriQBTsjAQqtRjPcgMWNSOo2Zk0H
MtvafdLem7ZflSYH5zirAnDuYYDTYnvgTGE1WO8AJZzMC3XcEn6zqNBpnHEJZunWXq6y0gehq/yx
GvdRQDxhtoPogtSJ9roa/L2q6Gt0vBPi1f8qRm/nBSQWzIC87Sb2zG8DACIeYs4lTDdNJnn3TOb1
K26M1gUe4OryW66rRmNwFoL6KUDFfJcn/4MHGBWKtFfl7Loo9m46lNS9QesH4yqZ38JCAGcYe4j7
3MX1g/qS4qK9MsQYUHUK53D+AzWwOrAhpHyIgsBZKgp1zvDDOPYDBjca+dXlNozIUxD7AOGNjMRF
N34qBxhaP9OSUJtu54Hpc11+SAQQXjfsnvPi5XvirGN7Pb396l+LZSrCqqUFx8cM3SDhk3Ck78jG
To7p2hnERBKVD5gKa+JzgmGmQpTdkSkfi9L7QVz4tsrgI81J2FTRpnzWY+tpu013IgV4D1mW4R2Z
3T8fAvnMvvzH7snIXm7cQNSzWhgGq7Y7D76SFNVVi2PA2gvXoWhkjH/1YS3HvNJnPwTEenZMqBMd
0MGkMy6iiqiiKJtV68RvJMTeU4oeqmfJwI8h4JoUeIHX2t043q02QxgfayXAa++aKFlN/TrRfzMd
bSEIPk56ZZuFpRoQ/OJ1zqZ4sCO4hE6vezn/v0P0+60Z6gnxqOIwTNUpgDQKKCUEG37d3LEUD9Rl
2++Qc9Nc79nD/uqktRulhv2Gw9h24UHSf9VICjuvh574rvaX+FEcpixrPerNO6X1bRn8k/n3RWRl
R3KYupwcZX/a1GGeRpHLgHQFm01OTKDjaSBcGbT7Gm0Ubw9YtdZh7iw23zOHRFj6L4wioVLO6CxC
vcWpQzq5tFvcp0gwZi7n4sA+OIraXuErcYjygJrQY/fw6utustj/o+D/dDQlGJPn7mIOTvcAwiJs
4dqh8we5AI8ByXxwXpbwvPysoSy+hDVsvoXQhpJgFaD0Uds8OdnZxqcqbbBDcZ5OTp1fKSjxg9dq
883yI5bv93xMECMvQkDvbeHv1d/sv8nZhfx5juMpSwnTt94Q2hE9XwCKrAzEsHVpij0ZAp1xWfBE
RoQ/vBiAYvTMBAaE23SxMCr8Vfx9vlEedEqVt33SUH24GejsgyLWMtWF7Mk5YAVOCcJh0fitqMsz
qIA3w2Pe7Mxr7tLt4lGkP9dItKiZmDyu0V20jl61eylh+eyabgZN6Voh9WeJP9qPHLJ+AdT5EnEv
vnl4ir+WGKK+cOKrUL4vlzyS1qwLkxUtlp0iroD94v7FfM9h9B4XMJmcDTJACe1T/IwQ4v0Ce2yN
XSvtahFimi1tJIXJup01ZHa8S8K7WMq5yxuR5JMXdHwObv9SrnpofPtLx8j5pStsDpOU+x1smflY
GDTktbwfFkd+eCKJZljhD4MGCFDdMtkhzbcYU1FWG9iQ8z2SEcDpUyI5adkBHwUGOs/W8N3auFAL
P6QZ3kN1+ZCaPEFaCQMfnPmftWWEalsNUNYFzfOMRgN03qE+aTEqKZKPUP1OCTPsz7Lix5OuXxty
8HZLMfEPLoxoA5Zhn+FZTgejObTbH44122CIF3Bk2ugAePGJjnMCKQSH521qQIHceMGhzdRWHE+l
xY2FFYtrxlUEElrfUxefjUgFJh99WrVokLCgAWvBmYN/WfrjzHLHKVWEhWuYaeatGn9rdaKpWE+T
zJyTDD21YnVd8Jsj2GoXoF7MN0JwM5USYo9R7YDesH4+7X9+7b5/cXUZqmA8RkheLi6DGvO2Plx2
7r9/JpVRmJGMzVYF32D7xUFqVQjK1pPUC/UnKbi+PqqxZM/PY7iF02eMpDdp/fjnHAuzhZaEH9JI
9L8pPKgTFop7FCFKsbsbXYicb6HpV0/mi+E+5e60z5Wk4gVQtS3HlD7EiGyOUUTvFkpvaAE12zBi
pi8euFn3ID95605SoSLSqJkVEe2QQffde/veyDKy07mbgl3RBvErEhe6rvE7kWTMP7pi5Y/e0Tga
uslhFYGAyvHJUX78QYDIzro5WxliqmvDk21D1OslXf4QLrZW4osPvMCOINJgzFj+7RrnniRSLbwB
JDjDMrMILeAFcEVrJEgD3wEWzNNWtTi5I4IiMG+mXM60cUlSLb8mpj4O5Rnp5MRJzmxOjdytS+Gl
Y3pgWZvEhGWtAXcr0D5kPyqx25wZUBgnC+eNG2q8NvL4CZftxKNeykMqjSypjb8nUtUxro1x7hI7
r4fCR74qwY1RUPTCxDKkpITq4GoL3JLZnZA21rJPPxtfuKGTPvW3vVXMOQ0e482l7XJhY84KgStj
vGPwRkHdeDEx6WKdMgOGHlUf+6Ny95E5RSFhJpL8kzB6+ipBDAM9aWJ7T8qWA4a3AFcq+Pn3sgLa
FTalZLkHHk7ude/KnjFALB/hMTZhfqTXci7rVKCUug9mR/q9V9a8bBtuRX5nVghsk8F01r0LC7eb
HmO73IiYyzFMsb6UACwJ1Lo1Nh1TuF0yt9IQ6CYqntGP6LDrgEvRs/t0WlzpW2GSCFz8JTkitb2t
SD9fWyE8nR/xPelYjztr+v2g7O3+jczbKd6f6ipm6hYko9UYljq3MRvc0Hm/Gvh3suDZwgiGo3Df
eRSoUwDskEX3lyPfR+/QuY1vOJ3YaQkXIXZ0WnNfGLH2aEOTH2/EqtXGGQRSpYIMJtgNVOHxeWct
ANg/ba7s+QC6ZHmGZeHl1kz2LzZd1oFmLc0JkXzAaKqN3qTvtcuo8LgXvHrmsSG69OCExRuzxjZn
WzejSQIUOHROwbM1QyMpf9v2zB7ylfoM4RLU1x3gCeGCTuMLqWLKH6oCtXmcM9JNsnWB0gKd85lc
Ib5RoGKpyRp2JUr6OurytdFgdhZp5o+JxPL2iyEdXZBGVeIN+YhUmJhigCJIQvW02PIq5op9tNwS
N7aY2F1oJ8KdigxWoLth9TF7fKo/FIrfVQpIst2PQVQE3z6mX1gGL0/T6YwU7SiBWIRgRZ3vJxAr
Pz5fTOoSDu3oqznDTeikvoVJ1Ld4UZtG5IwjuRZQU5eB5q2PSsmO+Ups16vlJUb6nHRwPxlgCsbb
uE9cOfu9u0mXPv0i7FJkKCZSGzYVS1m1vkhwDkcAl71UlPLQ61QCYkHPwsCYUD9ALJ18Ncg7XuWh
f8KZGi61fp27Qy27SZ5zLX0iNgwasFOQct3/Hn706oubrzEesZb8XOyk5DsgTuOhNSUBpR1w9XkK
RJukSQYtfpyownuOfASEaOv8MYH3DxTa+3VoVR0N4KSgH+JlP+8shD9P5gK2RoaxhpJj5OgMDFmh
YEH4ssCxB0zjvIicoIcmqx+5j9bBTkqC3ZQLARxLhvWDVRh/Lvt8GEtEKysy1v6JzR2gUnKjJm2J
hlmR5J9gn0+kX7a+FVtqGH9xdGXmsrBygV8YWfOI/IC7erGJPJtc1u2SoQs0flPN9uzbIN3QOKu8
GBRV1fQgdfALPu9K4poACN4np+Mf15NZ5NfkoHq70d66ugOus7uv6lOorGoGY5DENGmMAnbegJPl
dUmQieI/5wnreZKMhHzjddsfAuRBBLEu33X4EFKxTRGWmYLUVmB4LHYqTacDznTWWWFjv/ww8nw/
O8WRHoSYoI8i3oNFzwGQo5rqdQUsEqjGDp9bGpAha9oZmfO5rK/XrDkK3QWslZ3t5VozS33lQBkW
fNabjp+HN0b6pM290eirtjSkA84bKEuVX89seXYzsR/u8WpiJnXmh8LYkPHip0mApHQx/kZUOnqd
eaUbZIfk/3b+v2WSbfjuaTtOlqj4kR2vhcNlCI1mKkXcOqTEhg8G+9Z+r/Vzb2NciPM6zBmJiHmt
kazTTGkhXDu+asQrV06MD1hGDgSi07ELbblCixROq8ygASfEc5ZUEqHoyTH97A0y/g2YmuEVEWFb
OfSsvh3tyWejhD7YTJ3W1xsnwIZ5Nl6RYpH9gghrQxYY+YeEvMu+3iKPwv6x1zUywImTKv81aN+m
Mv7GBNUPieovkoEDwA0pDQBWPWuED6zAaAxN59pO8bfARe73KM8kkXRBQ0xsmrPRT1HpyRlIZi3A
PQU8A+AUfteln3KQ+Y/cCMnIxG8Ql9ZpGFtB3x87T4HLsDtAF9GmB83BqK4Fd4MMHpkkOUa2mCef
trL+qfBhOU0XNSf53utcMpCSSxYwMAmPi2LzBvng2Qxm5nq0cmEq07EIvSwFZJGq7pyI+ts6tqcf
in9e2bRMF0822cNixoCZSw7k6inrOvXsx33uAJMr2HYGCb314/SRZviAPW1OZmpMr/qrf7bm3M0T
pxnkNraJElqTyy43KQqMpiXXgGBtEeQKSt+SDydm/ikGSvr38MP54BUazgjBYGzL6QFleNIJBz6p
YzceP4DZiU4YMB56LKBgANodMKfWM6AR1TuCfUoNmR9lPlmougp4K2Vym8ussWzkJ3G8k1dx3FS8
P+/Jr0bgf5nmsIWg4VoZR8ylqyeE2Qux/HI6MKQ13c0pgfO6lXByxKWgnoUL0G9l6anOjgJ2LNUh
xD4H+/Suml1NoJY8L3Fovboau7XxqNyC42vIV72n0+/gfBlYS2Ehybc/u9NNECZMELUZvQTFSpNX
M31hrdO1oU7mBpu/nBXEmN1Z0Un04kHNar28Uw+hA+E6NyGnwH2N0qNqPh/92NiABVyYYeM5KwBV
99dcwpXCP76kW9Uc3XoiSXrEtsH5agCSK6nMz45rMbfRxIIvO2X1s1hcjMLVWNFsN00g6xMQDFYS
g7JA562dBC6p4bccoQieFcU9XMEYiwzwpgJUTGOjvo/5bWPslLdX1pr10Dr3WHG2QqQw+ve776Ty
SqWFR7kEa7ptRn7L96kdLECjr4vuB0tgxhNlsdNzsX4v9bbM7JdKVc9FIonzUIyubxPwwFKoKnX0
RHAlMRea7+fIzOlQo7QT4akhbIWpBup1dmks3st33YIrwbEf00DViHpZ7MVQ9fNTVWAgX3DHp08e
xmNRa45CroJucRkDYYR4gCm6tcOf4KRJRyESEufrVsqRQMik0FFMmnoartvALaJS2sg4Mc34SPdp
glWiK37+yCbkVvodgRay86+MkfUcGZxOTIFjAcfcsxwB3KFxVROggwDnHkSP0wU0yWfzBl2RRCv6
wTmUXNxNKeebHSYIXFKG4rIMzCW3YAlUKJ3Nf1j1zoIyiSif3+ZEeFz0UaTdISm7QbmhEVM7YO6A
qrzY537Y4Nm0BnT62KUQzOInSdF/ft2OOQHm1s3RKbT62zzjNsnjNVplWsi4POOkOWsirDlmTfAw
zwFQZgPeagbNeZkXz4x7zQLkmbbEhjP2PD0uQpCTi6Q58Gx3jOEqfetLt4HIaQAfME+xzix7sZAO
/dsHOliMtjlnUPu6kR9O/oKWAGAkpyU1ADIM8Scyar5MpJ9aaHvUV45IEm7SySkcXMpvGzk1nFha
3VXM3+YXcBpSkx7BiRqh0qVeIVfk4I3xaj6tjmvIKt31ISat3lt0BjUwptEWErHS6GcVLPsxfIru
vuEcls1zVbo3jnyfod7Iyq9B2K7TuphbiaZ4dkmMLC698RK2LaWskGxQfZonM721k8C0NTBi6qbr
euSXRRdVtF8yMl+KFG1DtOr3CIvVml/YC00Nv+D5tJegyluutDnycZtrtcwOF0IXfUHSSYs3n9Xc
54c5Zg92zxCBIZ5Jxyflyo4MK1QMkXgiiWOpsGYQ9TZ0kHFMfsj5yNvMbfi7A7PDBbX+dl6QkeG/
sSTUtuwfem7FShTWw1qoXekAWKnlmePuQbHuYYzaHAi+bU9dUumgQMlSEJV7lQqOZQfH3bllGhYV
Md2iP7y7qJ0ae6x4uuWA2DBSuBmhAJqDYb2riV+BxnB0lL44qF62mhjco1qxEB9p/xfwDi5Hh0ff
guhxrVaZrNbdupXDKsO4lKzI6j3mCkA/6anxwVxACV8burahaBjaEEJ+THxEj1bz4jaQH1MtYbWN
okIw1q4IArimNJO6GgtkoJPgvOpZMJFKURHKAX4YGgNHepH8FthQFfrLMrAweKjqbN7S1j3yxMeU
9PEoR2Wq46dEASMY4xSqE+ghHMCZKYcflxb1l1Yqj6HzPaoEI6DZw/BlZcSqZiyZpKsg5ctGT8sx
c6QHqVdcjqy+9r+a9mAoVspVZ8S2ArerVnvv5UR8MDFJ1lwZKwrl4fSSiytNT2ihU+LTsCfWag9u
3W6yVLcGIqAtiFkAkhIUSw0krem9X4g8K7wChy54nwIHWfwqEBhL5vQJuNKNOkR0CkxH+7ctNKTc
pn9r0nksPuVnugH34CPmha60WNf0BxcGwHR4JyrHRMMzKaAuXKpoNlLuAlwWTa9KOpjcIZ8yAAll
ocee8nnv9rL1mdvXvgVAuTc+YvaKXFIA/KmNwtylCtNdm7iwJ9lesk/7wtIoXM35YP7OTFUSQTyy
+jE428vOLd5rzveY/WfDlHlJ2i4IH0kSKWjDmWKqbloCr6V019vBz7cEaxseZXlf3/vTnstw5Uvx
hbtfAS59Mcvd1/If/zhxAZ9zjakUfwpDQAmDRAtJgqdD4rVtFQBQqkWnXN7E/fbzCMDgCIcjis9a
azA9qTbYRcFxnC2gG4nhZMP/7SbinUF4Nap8GKgGKkcjL+rg92Y9DF18xdGWR3gBSrva7WY9Jzfl
vHQoXu/zVN5Rqyb0edZY2rRZYEO45FVMS+atcylDBUGJHHqfey4yXTdiKY0bN3l9TyX5MWio3UO8
CbXULZJ/tf1ejy82Q/hcgLIupv+ZZ7d9tM07dmfVjQSM+TfBUtkn6ESlGIXOb3XreogZclsofwyT
ZpSEBlCXSxMNjeQmM+m7wfjjUNKfLqduqQChf0hHIztsxkqFMEpO+5h57ndZzxivegvVfMk5/mdm
j7yTAYdtVX2HWYm6TjoEOcvzeBT+rsq0xY/CCoYMaGHvP5y142aNAaF9z2n1iUSoqsAS1EAifnUn
fk91OUTIekRV1x5pFrpNWGOCOwWjtcO5mOtzS86/xbA32FlcL6suMCWKF+iJUJdLZhKvhcidfkZM
3CXlCMzgc2WyWP0Oy8geb1tqBQqgFeVMM4SQepgHuHOtdtSt6MweAI/EtzRTH7T9ghzqTfNFSVAM
hfFBJARa3Ke8J3krbHdXwVMPNphoILtomhdie7Q15yF1UAbgcec6JIpe9UEoof1NsHOvSUSekfLI
V9dyeleNRj3AB/X5psCeyrI7UdG0yFGumsybrG9I/FccQTsLjg3Bpdll0ADW1FvhULiWJdfcIgzz
E4J9oUncFy1F2NKEzwQ4wwFQRRWKmstv5IMTXSxF14cxloup+dhG9UzTMlp0g2knwrFeNKnK357p
ym1Kng3DRv/bkuHt7vHrcqpAhihWsino9efBqCYUSDU3SaOGDuUoFN34aS0dbyrFXWVlEEMM8Vbx
Ppks7oznM4hJRN+RUq/UKC98MWkBz0CCYI3l2bZN+RIOUdjAQAdD73jkFpXxTQ4ZUKI8dNYDWeN4
UUcLkZZZozs7RaFtZ0oUJKeeJFpEqQe6LqjgtoA49ktGEtsIhbjoFqwp8f9PHc8BOiFbT6sg2YNN
Nl725KsczHz1iTN0gMuv0UHuufztJyrv5FMbSTVc8opumiyHVYXG0m8Ibvo4LSUijgeEVM4Kb385
tucW542NW+Id9PyeRvqXf9D1u2d6WevgDCmQUuREOfjYsZvJweHxDw19NHwaIDt3LQiB73zj/ysT
4tzsEoihjGT7bhEnQbfp2dqfdsR9yDsr2ruQXlgcphXVWq5I2ls8k1iUtt/S8Kkc9T+3EsXocziw
BvSgBiy9THBW1w/ykT/ELSrXu17yd/+zvGUFIc9KVACz9NBE+o4QuUhpfqk0J6QvcSYvDXIWqiJc
WytFsVk1HBhBTIVIzf9YC2KSaVSAe7073hlJ1XpYvobmmDj4obJqAltZEaew0zbzZpwPQZ+oTE0D
o0dxlLTv2GaMrgQceAPAgDr064n5n/z6nW7FozhcEa/+mwZam4xkGOlo/wW7nZjKWTVpi7fhOJxZ
GrUwk2H7l95L9kbj+0dRNLjKYwiYRSqy/hGISOCjLf3kzhjNREQbv+h/DLUqlnMht8E5eRjGRAjM
9+ADRotELAPFJfqqVw/NIcgKlEiIJPyQsy/bt58WwWcfDoMpXRqombvYzvcJtvpw5B7icbEypzr1
53kCtjJuwVKlW1Grt7DKS0Rxql92VJ1br/qVEi6EGQmq8VpoVAWp0WSjis94oKXCQQdPei/Ay9aB
EjwrbLxEQbX2CJER0t9vjlwucpDPVanq+RlJKxB+C82O59rW7EpqaPr45RdHpMUJbexZPK+cEFbq
PTeRgV2hOjq/3WkLEQSizzpVHw7PPX+n40vKCNs4C+KKiU8lIc1ncZ1GtqOJX+he0C/SSClQ5cjX
ZwhnauRF2+ZKpYMhuMDXhnYIJ1Ytp5PGUghTp5rcU3nXREAcm+3krTvlyW+vyBmsaECNjvdgyeq/
uk070yHytvzzuJQy79lHF3CYdtFc79pI6XnXq3yk3/Dk/LnhhGIWGjn3oQQyjNzFtbb/BVWARvpL
vweJYPaxy/HCLl2osHDG8FBt6W8gCqsbl4874OudUvULla3393elZGIIY2Ltf8qSRYtzDEl2gKFS
l5/8P2/nhuQLlQLrBi225SKlYvHzOoxlYELqc+aUuXbREE0h7Og3Lzzha8l+ovxc98bRpdYqZdoM
xooa9UdEDJLxQBvl7rM1y1qC4zj9NuAEGsJF7xscbXzDZ7KndaHcKdHv7+56tdT3iri76BF13ZYx
al6I5WWMIJG9fPKS+NQ0GMAnXj1XZ/Ya4omzNES5GeHuzNL25hl7BIkgBWnQiIoVlpj5iUfMtCw7
XMJxFDIl1FZ2gu2PD1PQIEDjsO68DkKhzNfZi8NxSIGRA1GmZd14vLgNb6ND+RFnSJiyWmQ/tfud
B6Z9KQrgAawaxxdzNCsO/AqMtVmvquHj5j9NDWK/LW5WcCT0BaNwE92v7kbteekpJJXcAqaFtNyr
NI3XAe4IpFBGSaba1hIyFSHQFuhWENGvgph17FyJfUPS8AaYJjH0vOh6DUe1xGI0gGNqPAZ55Bf/
Fl9GZjmruSbNjtYhiGShCGejHZALJEQ5YBr1vobkhNe6dX8NvA8Z+KASQqt+2Uwbky/sOgJGaR0b
YrShpPpkWNZuNokNgQNo2KDeMMj8UPO3pjCyJLHfxVP18BWCsMYC5QPXsvDso7H2R1JlwDkapxny
wJx9C+Yy3sD+44L/qWDdu6olIYhfs0xzrxzFdtriWUcWyXUCL70NhNdrdMgyvKxYcaiScjlhNm0A
3aYtmYpRjkG1Zfo1eA48AZ9aD67tXhQQMSb9RHBKKNva64HkT6Uqbf7WpH4q6kAqsfnjG/WOIQST
LrLvcy/37hFXssYUJtj91ktWhdtk7zPIrxKUi9rb+B8brt1FOR5odCTEIW540UO+kHDIM2J24zqF
MhGsLnwd0hCyQxtAxx4EXOD3EmV31YFknvDsFxYm2IUesOFRvXP9PkWGkOTo6R/YY1hsFNO+83PB
0uFXBxJndztlhqv7DLWZGPkO7fghD7q8ITAdIAjMuGJVOmCLYBHBBG8OWPBtONFI4pB9VvxedIVL
VKpMgVmNQqpqHLdMriFxvaQN1+/xUBxy2NvB5mtYWzbIVBUULWnG9PK5KEWXBy2BJhLIaKXf6dhp
jHfTTYErqzHERQuJ5VGrJItcVA/DLJ4jSPUoqlR3NK3/nnEa/c01V0qMyYjpybdMDNG1eCu4CUw4
aimGsrxRnPxMwptNGSZ902zAJZzvFq/uQaYVj1ZDOrNz+mGphvm7sy9rrzL4plQet/CWwQTF1YSW
AdEI9Kx2z579fTp7rE/7wY3LE6b5iXD/c8U1+q8sbT2kLFWD8J+BKFY0cc9kDYlk2G8dx4Nnbz+8
UJZHilQz5ksFaitVCJGE270V9DCjNH482jMDUHyTr+7ct81CJoYDxyNTASfsqqezdgTzZnF1MGLu
vhDdwcO22ZgRwle+p4V/48wp95/OULpgmtp47QKHbmRsN6eAUkFD7nUN7ovh2kN4ltq7UQB4eJKK
Kr+/PlnICBGo64RCDh7Uk7u/VedA08eBH3BSACdH0a0HHG4hD3lkHF0Vr/tIizOhRp61ZMYcRUTZ
cNgrwzwWRPNOOijnTcuRmWp92kivAru4Am7VH6V7hAmuSoTMMQqV9zS/NBBNDxxv9/GecewVvjVn
d3G40vl2t6YwV3LjKzhhJQHxnvHOykDqxEvLXaHu5z0jSj+u6iwjeXdJLbywYhmEstyd0a192XQZ
CcUb9HW7LIWDNab0P4UcJH5UJ2e/zWyk1UFqYwzv7jmCKNyVoS/row7UCQuLCro2xIXJXqO4lJ+J
ondTL86D84LWmODCTaBFdUSqwqp/wIkTThr6kaN+MmMW6SOXN8hyBRj4+AG7CcJ7f7AOZZwULG/s
Vwtcr7OxqFAzFNu5KrUegNBvnBJLmDi6uhMGBC94juQmLqwtit6+yBCaq38JK1LpEPXa8FmSv4NN
Sib7Zk029YVO2y8jj6rZXueRaEyuOwYoSSAQe2bXsb4JEiFlrBU2OPEWG7jp84V+LC4eK+XTmal9
vQCJtsPm6l/M5CgZODnRD6atJHTgnTCK0zYSIcMe0mnjJon/uaI76oAUhcZX7EgfXDogZ0U7XgUA
f6wbnZ/SPybskRAg9zSMquXUHo0LoDw2I32er2nQ/zWj1BEy2frbaJaS+LbX9TiRYXKrM3Yh6zNl
of2KqLJREDADj5dp58fK0BVxlNMk1Oig9gqp7DPgn2ar3NMhNh8gTbjiyWftTIIlkZNsaSBNL1xA
xCDdQF+KGUy8adSDRs5b9KBn4AstPd9NfnL9wgU2UROPb01Y2kocYIQWR6MRf0FEKNqdamRaLwUv
Yce1hbcoMk4WRRk2TI0L9i3w6BdpBLHpJwKa1uHm3rxAsUzJrbTnIIYEyshIAuCoxGcjwi+uiyOY
zW6MtNq6wMC0AKFuZ3ryQeyi1f1v+oIW7quV4uTk79hw3CP9rPEsIUyNaU9ZSIyfGrAi3gX2DYIo
v2ggxLrMYHA8EK/ROUIrRqEZa2LoqHJ1eO9J2iwEznjSYCZ2kBp2gBoQHlIIzDFhM6HhoL3/KS8H
D02JiefGVARUq6kjDV/BkBI/KTDTKbuFLkUPGsb8mfT8aMDpHVM0eLjdZtRTkqwlzdXU+wOLkKSU
FXFzVKMZYxR8W1s36SD2YjfKccmrtFIQ8FiCeILtVVxhCL82YT3idnrIk5VFAE0qO9/MMWsn3Q2X
guJXIDMZlRAIW0q3pz6KSph4wp3H4xu+o0G0G9jvqJOuHNQvnGzhCQUY85nEV6qnkssZHO157/nU
+30NtJWdFvoXlIbH5jVmhv3JHSooFEaJbxcMeiJ1VKxyBuNmQhQ1hnAxUgQjZFsFODoorfR3TV+z
O8VMoLgUXeptD14qJTGif6r1JPwk7nVRMgWDD216p2kBI6RMeacgaVV2XQzbJwMyX8/dMgBqq7Yx
61KU8b+he5lIrNXvB/K3VZ027vXalkmC06LSC3pYJsUprOqURcasXr4gabXKuIU4P/WZmBnztnHw
TjzrqQETWg+Z6A3FQHyKSaDyaHbv8/7YrE8kogMsWhbMCgNhoPQrxzBJRWi1A52gpXLo1piPOojW
q5yp0xdeNv8olfa/cWBZwkguHOgAd/JwJNLNS6wdaC/FOte2TWZtyaOEyBOEHLAiT/ygr7NIBzRr
O1nEgYk65FjMRR+nZnDtIeFNFKwjscN72adU5kTgMTfWVKQ3FOZXdh+mnYHWYDaWbfJt9w7XGAmC
j0zr4zQEeV4plbp7cElH59eFNt1uHvhGwTiJVfDQPXFsR3FZcEEsL7VcGIlIjub/mgFWxtnMwY0W
kYVz5VZfhnwkcfKTJnuIcAfFbud1tQ8iAcQoYYZA0EoSOiDJyi0WqRGaN8P9Vfghdv8TUxAeeVNO
rXXlXwxwFvd/QYvRLVB/tm/T3ARW2kYdywouY1hFAEDgqmbz+K1z2ZCPFaK088+lF/pxIdjEi3HW
/IjjJD3K2+IAypGbamftkMb2BXclgjBo5c284/6WriS+4HioNR0X8ADF4mkqGouOD39AQKcbc0qs
ijp61HqPROQ8R2BbUVtjwaSR3jJOf6cY3sJpoFKe4FG3eQvTg1TcOOW1alY0sywykDcrO/od/fDf
zzF+jAfXFm9xWsT1+X+jBIP58RCkAAAtNZHgO72cS0VzvjTPz5OSDX0nhjZXeAQ4gjc+PpImttoZ
5I2cbK8vhGptOfZrPyH3TjN1cR8sf8kTS4ZAZRkzwzBzUVDSUMKHTnGUqahNyiRE6ny02YfVp/ee
yalks7jM2dShBDR2TC77iNN1EL1WqU8cV1Hb/Jwhphg6VtIrnGbDLJzpft7U2Nx1plCyA4vFjFnC
dRbXR6juqx9uJTnPK05zGuYehJN0Ww7hKLAtViZRj0D0G0YuT36i64E5gPoV+XyarlTPV3O96dxs
wucKcMG5ci2A/wmgpCibQpua3xqur8mV2ZrqK3+M4CpYqVnuipmoGwSgXy9Q0lZ0fXZAxakqRh1l
NhL+2TMOZMKtY9yuDFEar55AiomBdUbZCU0v0B4ySYERCzZ2hiGQmZBEuPvjTnhYlRZJKgjqfIt5
iTx3BOSbTI//BMvCzIcfoUqUVtmYEJivUyQK4e1boFM1/G4BjQtKoQFYY2qyjAATU4MhAKX56wez
hgvHVJWXDyWfVpOoZEwOOGmEP/0zJK4dz//uSmny3IxWmGvoo3rSb8Vk7fzgx52WJxiuj+Hlubvi
fsuhhYsZnLbx9dkgpypNo7W82bv6BJErn4l8pxjLSHLufTktYub2bfK8sQnF12KUV+ywYpU2XXME
/LxDiYj09efxW2ANy0eZk1zz7puuUfpTO8O63NrdVnKQjfhRVnTD1a/aVAJgla2t3Tp4TmkWavPG
zTWTcbNj1mAY9Xbi8kTcI6V2AoYqGAs+KRxWcxa6irfDKue3dMz1Y0M2ax9G6N9A8lFVErGkmNPY
jcdjZkMCrNVeX3h50eKSza4xSmHTTUYzDQFGcCTdEdj3pQttrVIQeRFLCSwy56TJ0TP1BoG4VxnM
pFEg8lauIQIvShS4T//L8IfifWJMFgF/YxtgjcyUxdm8CRcsQ53ESMrhRHkfItLjc/iqMw/5EwVL
EaHo3SC2Uwp1bjdPW/UFV5Do0LFkuTMISMfXMJ8U/Zl7i1B/1zikCZBbGmQO5cUeGiZfPbazHA1Q
lMZh2ELc/b4s+T9bjaN1kdljXNWoW1x0dtaqB+q/QdNaXwcpwFwUcmdRNVHowLWGHfy6xJaBKSAc
ZHQ7SQ1G3IFc3xpro1eZGq5X/dbwre7obJcjr+hDU5pnb00UIbeMQ5kLqPtE5oUc6lSQU2oeskE9
DAMeel9Y3jXzd1C87hS4TkTCGUFME12cpn8bXpRDzY3mOnt1sgII6Ajiln0tEF407CJB/hwTfMqk
tjjQF1yhcoW7qLFG8FVglCrippiG+sVrOjWByXAFrnyENfkKxp31v9rdLkE0+6/tk9M1Kp0gBOe2
qATN/uaodgjs6cGhB0nnDExxMeIY2ymWwElvPCWt5VPzZyu9S4NPhn1sbKFGM3jGLrSOwvwTSrZd
SCy2ao3SFvaRf6gVPyOlaK84WqOaAFy1u/KebDsrAEr8YxW6IW6pvmRolamhNS5uWIVCFpsTiPuv
x/FRDtT+1gq+AgA43o9cVusKN0O4iz0B29SFGu1ztvM89gaZ9FFngz//FraUbH4ljc47vWSBSozn
chD8Nxq+Aw4w0W2vWNm/8sajKZwhE1Yj1Qmad/mc5s4ib1xFVSBnkzc/Ohi/UvwKocZcGdgt5oR+
EmD0FBdg+bx5CJzD6caiVt9a4Ma9eOn7sZFdwDQe3SgWr1F3/Urps7PUlxMvc/IY5uwrwLV9SAXi
T84i4Y4x89HnmGNE8bkKZFPyyb7I5oIbix1EpEhQKjpgWkus3LvS1pdTOouzl5LmcBNBBTXLMI47
Cw09zphK9niJ9bIAv1f/SnrKIcrr8rw+ZiE4cNIhWRi9yJqhdupelUE4pfTbcjz+3JmzTUq/VLZu
jj16K9F6Pi8z9/23t/GfABUWtZl187JTLE4X+dVhxnGDpWjlSfyyoCycBBYi1JDz8tDhWtGz5BNI
IxWXt/BLRLPILyyWb37MpTVX5zIj7ytaaMw5a697S6HmEOC1LDXHD953SojW9pfndIyRVYzyuh8X
9z5Kw/RXmGjP4jAPN7pPUvUgq7vMfGE5ZMJYSe30OQDPCKPD0A94aFHqLJa8es63ertW2wlqnJwS
7FlH//HNNUQxvyEUiyk95KYXJ49xMg+XH2SaYCLR1Y5MBqbmhJhJ2PD0uwXrMyD5BOUMNsivtIdZ
S8g+so7Eq4eGgH7DjeHAu7vGN6LfmzfXPaSI/QMXh9U8C+Px3CQH1Yr169hdxKiOirmIWbpL2o+j
PT03AkNFod2d04xxre9CotBPzp3vjpoM/WCABz5EepWFlx+BBb9zxzA0BA8EJQC3DCl4BqIigxUs
g1yFjsEi3quvZr01h405/b1t6OQyQLXgKKFxNew2GLo6KVtTz4K3ZieGP3vylz1m+BF65t4EwORu
fss2Was/ubNi7zvZSp/qf8CeLUqasucxT88Bx4+Tsrg9k9n0unQBJ8nBjQzWP+jrtYHJWxCmGL9B
xOEnNlH1e2kmFdpHPqsNHGqSuahPF61G8lY/Azz6u9quCagWZQ46UPKSwSmDoGy0+nA5x1zXXPS6
+1T96MpytcdIMHVLZdUtFxE7BYjHqZzdHOVWmSpwGuDGPvRGtfrsvGwAY7mBlEcNdU4/6+sN/5yI
Q0rDsHQQkZQTV8MW+H3mcPzQCgwwzYPT2w8VNkPIZRLFBvqu1XZI9O8wtUiz9ZAe5mJ85y8TjTj4
vWvfzwgslbxbyzdZ1t82FMw7l5JFAJwT8pQgnqn3O0262Z5/3X+ISdlsJ51idRNq/M1Tb06TYOc/
nMsN51IqDyQZPC7d/Ary7PG9FveA00L9gw6LuyyMjtkBEd57E0mMcovcuxS2D84uieXHQQ4pVlbr
zrbcLZUVJ0wCSwlW2xLajwZrebA79gCCHQqt+uqsJqTM6h7sc5WkHE2Knia5KMmzWI0XMQWnX76M
D7+odOsXXD5L/zB5Pnjj1C81GcHqOM7BLjhZppZSy6OYFMEC/R6DW8Dl1014K8w0Q43/nOI42fzU
GrlJq4GXeFwxWaaRXb4KdsD0UFv8mTCwDYKBcG+jJV76/EsPa3OL6l1pi7iAVn2yStd9hntqSm3p
cEtpeop8Rvh+TR2Z/sOCH4wuB7aeR4HnsxOzG6fnMHFCMzrtSks1ICWgeepRMZ1ylsh0fbWJ4JHM
LIgcYLQmGVRBMMw4VOiFBCUaGUDOMlqk9xajBRsSliER6uN8pKWQRDJ6JYYTlKbfcPjoyqCGBItC
pb4lt7ikxb6FAvT+KucwGV6RJxLo7lbTidXp2BcySUPbTEYl0ArSD176bU8Iya/wUHWcFCnkTEFp
8Q3AaEwLBoy/di1SIF+u1nU2ITQJudZOKrbKKD29MfWjuWaQzjm4IkrPnwHQCYyx/itbvG9kClOq
LM+Zt4wcs6hGrBY0kRMPJidN/ermey8kzYDmPXqoO5vmvt3ywFkQTTokZotgsExqT5O5TzT+MgBz
SGvTybdl/it3zC3+dsRviMf1K2530qPB4PZcGFo6HqJO7IRgy8EfgFlb1x237pJcao3jeGj6aPre
ouzzFGi2Fj70r3pthuJp6oK/mLy4rQ+PBTlY449RjpwWYj6EWj/S8Q9kCBHGtNDzjWNShObMfxSU
3VMvT3mNm4b4Ff0/NzPfCEZ0AQMehtmx/tgzJlmtx2q6BmkZZkc0eQssK5jRQN9feCd43Fs6hiiq
4QcPF9BVYdLID9OSRWH/FF2trMCzql9Dk1ELQHkkm400PjUjR/0TpkPGcLyGyLRsJMNU3iv9soiM
aDhc1lwrNRT88ALMDgH6eTUyYm5efebJZuUbjde/Cwet/AMyIYEPIA2iryj6z5pmy7hXIf0Y+cXv
/z1WBZu0Q+TRv0JowwdvA2SnVbnCKAzEINBHEmHHAj90C0KVV2ultw5uAl7wbAX79CKBjlzv3/Rv
CRy4rvdh5e6W+QOt0dqkuUbL63geSUpuJtI0W2F4NUny+IOscrmFK4ArTqwLdQJBp1xVr9nuogSh
pPESHPLqXdqVx0trxA2wHs7RtEr7+FpTnyNP+Caq2ft88cAejysxfotUXfpMvd2+8grYsokx/SIE
pdh1wDVKJWmjvj2gBU5LarqZtlKHjiChesMD4fj2e77BhrT+GJdBADsbj5wCwlruKh61YGn1Km9i
VhneD1M/glB5v/iiMGmWiO9liezDoLXrleuYAf6mRG+xcxcYERMkvxqVTJcliDvDdpEcXy12NwpU
F75JU1s/98G3GafpaW7FLNr/LsGS+FZTegedupjvxQKxRCZG6A7zGJYk2w/andSJ6DVGYdDavtyY
LRnjvLtNWNJtr3WifdYJ5hGOllBMf6LvTGdReK4Ngl5pdOpfA4aaHFwVRXZ11O/NKJxaKBLmM7EG
raAk3oNsx9UfFZwC47SXuiMauAXiu8YVekZoIxdTiuTn5tmNGp14td140sDPCp3MpW19yDUhkgGH
rBSyqpQyQO69exkOmzORTq7LrrjoeIyJnO7BsRnxN0+MKP/e6rVT5sDWBXn280kmEAoxGG3sql27
yUYDfBEhUfsGn457YcYNU0Cyyzwi2Q0wWf/UREcGgTGb1iVQ09wZf0qnRZnjrV9ieaSKzCbqunja
7Jf62KngzT6rLtOTjdJ+0Q6apL5+c0uAsbJZPLwvreCknI+TELfvxArHEYhPbQ3b6JCWg/K24Syz
cg2ZtBvklk67pak0s2NudMq8VqptWTcIilfYBlRJ4phHANfHhV38HUP53XH68C6bMUAumdDsqGv1
uydob660yu1OZyIFhv8nX2k2uz8pI2hhFZJpCHnTzwLiOwWbbyN4NgVUjHWApumh4GZloO8AFmtS
8smTAXYmZoPkKvl0OrJa5yU/BzLIFCcwMnlsHqCFRWyTVpJOHBBfrlL4kBhmkfd2As0AoO0NkFBD
VH01sX1Deh0u2sIllLlOmeX+1u7xRfbtSjEEcBGMH6wiyq3duyGiqqdm1/ZFkgZYpDGMJfP3gd2P
KZY8vUZHJICULhGck2/X5cMtxe6SVzVjRV8HRM/ZYzjotKQASIHmWFjZiUmXSecMotmLK1s0Kj+f
viAWEcKvpioT4kDZy4NxO+UwedUiMm1AfQCCNZdJMHe/LLVNNSTsf2On1ZP/UOfL5kiG8vN/laff
JbrVDDt9vTS5YKmNfH09OGmLB3caFEPqEtIe6FkyyMv+wcQ/CeH9uPz4znw69eqJeDqz7FMuHKZa
YWoegcvJQ3Nxlr/wZoW9Kwomi+TUMjnCz0w3WnNsk4b68Q/9x/0T2hNMQLzi7QMEcCACDSvjAnY3
M25v3g5eFv/R9qFJPB5ENnyLhlzfEFIgQCpCGB8MoCz3JKsg3pYi8nr3LW8LWkKmIwlRsNaFf9bi
DL1yw3ECZ3HcX0662V+PuOaGSgPeJbEtfBSMKz8+3fPZwua3HOMq1Yhf5msTXqXJSHrpe1pgn9/e
klE1/gngHKnycRVNUK5rjz5YJWT2KuGu7EMhOxLU124Fo2WJEg/ePfovAf1jXS6E9E5LLFxmh6pz
dwO/MyjS7SsiuZB3B45G5qU7ZWTPMbwYhzc5fjuonscFyD/HMWM2zDgrztV+dSggMQpS2QflVhR3
ScEVJ1msLzajal1ZVC4dDlIt1GzrNYeWp9AsnAoRbe6XbGFHaZZEXtrq3DiWYdZthW1RGQPK3rrW
0ceqM7j4yq6W2U8h/4N6lVo+/k3ylogwzyStRq2QIjzrAM4ug8RrVNMLkshOQd4EnxCLyPVyF7cv
LKJZgayjII7H6dF1N26JCv/7uaR8zzrs3MXnMHcxkbAf2a7du8wp6mmeFfd7vqorRETiq+2WUQqN
bcGYCKaVduKAz4tQiYlgGC00GlnWW5/eHj646di/QGjKrnT0yIkcDi4MH2Mn4eMqXWQ6KPX5XKJm
zU1Aj7G8mYPIQrOdNWy5m2zRYDnjKD/nGp4ybG4hy0dU2+FMn5khzDuizv9aIvI86Q7v8c4QjHv2
JG8hcHcDyb2IQmEfWqTKsgqA+V8Y36xN0lBn3BdJTgQINxaMfhXL9AnL7ue+Lke+mLKyviuJuQP3
yb4NlTX1D7RqCnEYqp/bu6KfTc/w3NCYC8eBUDLKTgo2DEuyN6k17kjvaMWXlO49uhY2FfsZyiQD
tRtFT6NRjWkeQypnRw8s9DwNmnd2V2CfnQC8b8wd0H/xH6y4buOkTAEJ/xNCnTFPrd3aAFlV9nwP
TjEe20nI9CFXI1s6QeK2YSuel4DsfSOfwWPuLnUEljIa8mexSD/u59fZ3VIaWrrwmUV5xrFOjgz7
N1wTJwILHpQacRomSxQfRgvj8WtzH2q2YY+60qm6gnRMY+BOgRNPXwUlzbmPEZf/6ZVaAF/xn5WJ
A1ydYVPATP62KFFNPin8PS2kPiTptykBuDe56PDhgA2ezc3liMr/wjqDa1eYc192BDuh65XhIVTA
X32XPdCQ1pRa8Bi2BMzUJfLveRg5Yg+vbl1RxjiqtpsWrfbzM/VLh+Pn/J6b64RoMJHNuO7BqWoH
VFjA05xw1LbZPoYWYE5mx+8rX449ATiOfYA4/Hu37/I2CB6behm1fuV6daO+qcjs9wFQkkPx7JEg
Di5UB/MevlOKq9sgnfrompYOBA9HD9TC00pISlekUnsQvudnWJkvARySLqPLQyKtg91khRJPgOEa
mfTzS4iGD7cpdtZODJXvlC1aj1o8/GHQOGT0ACBWrW/oYHWbDM2qUP/q4WfjNBczR3HlP/Q9lqL7
zDBHHIN6dVxFLCuWzcxms1xSPwN+b1IiTKxBejGzkWeVgw/aNetJ5/8Mfw+O5DBxEkI1fGljv48C
RErT+lMVQ+wV5syXbTHGesTUiEjpeeguH9zxLoWSvHnssGyXmYyYNa6JMqkPnSo69tp7a/cBGCg6
EXNMxZfobcGbmLI2hSkAhfraHeeeNgdOKrzMnSFq/NvXkDuUzKv9tagooG2g4pzZy76EE9WYe66/
HBrl8KEuhKKX8LrdoHWJhGTx94tE+KiPJS/1AVAFqyVBZYjCAWLXzT89PTOB4KjKbesiMtEdWsTI
eRFZ8CR4qhEw+3ol+dkIiIPXGE0Fwt0E9ZLDn6M7UKw+xOUTuanbUhn5FiO2WYRdnB5g2bzKiAY3
DwsWFnaa80QzQ9BtIV1poV49htXHRrsZp72/09TXpqqq5uxj8aGfU9GPi3sF9JPOQaRqhCWiwsT1
kj3OOT9EBkfTy7Gip0akWouYBs1F12SmakxGfrRYkYohyxJ0OIWNnfnrU+OEzTMkkil3ValaxxHl
ARLD5fXW7umywv1xfqeryE8e5SZPdRD2nO5uR9h4xOztSJrnNu9f9alk1Nu6xOp2nUMUEuudyNLI
9sVPD0QoPNn0eftnyZcJ12L3dopnhCgsq7WbtaJXZjmGMpZFSa4zAkpm+inJHA+ZoeFIBeVdURKD
SoAAasTNtC9AfQ4gK3Gh6nyj8LIs097STiNwtV7XvFO4BvPanbsI2eYXI1pBnF+j6jHsQrsEPE6r
JOOPGPyKDynExSBd/5yOumzWV4Pv3GspuTXWBjiYxgdKyc+aR8GgyULeSzlu7UVFPOOwhaG5mARB
38ntVlbBRRnqNucd3maWEw/XWo42CKGSgC3k+xr21WFri9EGs/opuOTbru+GH0hNSwZC2zokHhHo
Tih0B3sY5jX23D/I8v3EX9YpCMVG8HXh7bmLcwSxujkZ3gQFNekZ+mI6BryoM7NqlyeRSJMT/4/r
29hYmjf8zxl5ImDh30dja0jiKRPRPijGO4+RqgBwu5pC8yrHwqo1vlisx1855y9FbcAaUlDXVK8/
m5qT8ipCGhOBc8MdXJWDCqkzesKBjq2pib3YQ/D0/hhoeIA/Nw+LrCfj1i4e5MjpBWv9nGkHQsjf
IWNoU3F4Tl3kNv+o4RIe5Hz6X35k4YZ4kkRkDeRtMMNEl/NI4c8MPSqBH6Hu0BTAJEbRm1GwPl7b
BpDxu3jTVrh7uZSaW+Aat6Gx5kQwiOnfnYku2gSAaWn/2WG4wBYS7DuqfirSNarkpyim04Qj04ue
r5M43xfdzRMMQATzNtsPwyE+zwhQ5xCaLHCfvdEcq0AIm1Sn0h4Y1lhSt9ba8jGh/IqnfB+PyGPV
CMP8cS2RrQrKDed1fHCw8gn6812dW831No3u5ueDzPAQxRF5d4yo7YnpmvyJ7krvLATSp2ELvum7
3LCP2HQsTFE3y6pXqacatuBqjT7BCaRqTc1qdMKA7gLBg12xMi6FDHbcTWoIMikVihR4phgROHsE
OfpF+auL2iYndzDsehYxvON5ObLu7VdSboTolS3UYOotoKzTMOxQuqhyVx5U03XJ0Zc7CxBRH7Au
UpzqBEU6ieqFUzQjzNc9sZW/qfu/I+VxPvWPZpehs0tHlE5thkr/+wNXw/SR/wZ7i/Rq+iJbRdsY
gXBDCLch5B1yhL3cMjUTU22u8EzL8SEQQPlUXPVr+mkyssDMoFyioNYd3HoBHwlOPMm4Ge1XvCOo
clGmRpPia9hsgoVSOuJ2Nq8HBSBcenp9KqZrBsXhP6r8GDWUOm0I9tuzeFE7kQNjeFepNowMARmf
rBCen8WNtBKBo1BouJF54D95A2fgsOtB0EzW565m8ABe+VuxiVgpJojPFMUHybvZF0Fuhc0K67Y1
xdK4GJKSAK+MFYCBHbQ8chEoC0vCSqKtSvG9wPLLANwCh16bpWPfUdsywfI0862sc7LrO6dfx5bT
gmILLldyECssbMMrXAJvIjTYWe5GctAWX0FYY7ZUI1FpriIEMc+PpK0ukms8NnF82uSb0FEW26Q/
fozQ1AcDDZ0y7llwFGEMyIgv81FCN7BL60+yqA0kQFXjImvb9oEYxdSMX2m0ifmefonSO3ZiV3vn
e5yZ4d/jhtxpbGFUev2HAeI9j5ISmQvPMRtVPIJj8b6/SZOY3unUCz31ovoEl1KU0tWEkFG2rv1R
MQLI2gsY5POByCNSKKvXUVMJGN3i0SurDlkUHdYxcwzlp49jSKkByVO9tZhjEhqbmfTseGUE0RqJ
wUf+oKWSJ8fJnYqy1hgd28aUEVeCm6qd7uSYOTrVnQj7tkkLFNOmeAiXoYfINTOh08sRpe2IflCE
uc5+mst2xkWaovfYhV00FNCM0RGEqxdCPE6ScTP1NfDd9dnGzk4nuzZ4ixYfO5C2tfneMja7phxt
YXQsWnl1qZNAR6fQnfW3b2inQJPeq3F39Pp1iCJe79s+dTLNiPS/wO0qJk6GyqIJcq8LErWXfAcC
jKbLEbBgDutv5TbEEzOj8mHeOtlPpnuw5H/jOO7yDZ+1Cnb56djHf8BvU2ZLgpfjza7RlXtkoO3l
e1b8SLfJREFx6ojjuqV5e3K/0IFokGixNrNc/1qqJJ7cAnOid5ea48Eh7Qzp9dr22tYoihFuAcrH
rHkw33F5GD6w2npikJHsMgk24FUN6Qv2QI0+iwVpgv202elllUkq5CUf/OvhmwlS0beBLorIqLfQ
tWaMKWMINCZbbr8E2jnWI/2JN5PIlTa4vUBXA6z4yc37shljHjGKXvuKiXjDOVDoQIaB8Ml9Nla4
cayuwVuH757v3xc8CC+vA6Tq5dx5SZk9NekRATxIHKUwtKGc6oQAnbJjA6f3cVkBaJ3itPUYliJx
Ys2EMSKSCtOu8MDdwQINDpnpkzY1MYHTImytJfNdkB5GWK3kg1f2BD/rmTq3YMNYSG9Oetl0qY2N
r/RmVdnxECAajvyj5Vrsr8H6mJzbZIyAzUvdnM+2uM7OxdCWF711Z9plKJYpYw9UCcFSptCaXHJj
ieDVwPJ4ZbiIpuHz6FmSvA8Fn2HDUFALaP3mp3eZnaaJLwvOxkMDrQswqoIt6cwJBMbfiV05Seg6
GZ+tqC6bXaNkBOnL6aPYMFueXuAelzqFf9hwMJgxI9T9ImJNtUJiZlLwbDscpuVTcLMpqZ/aSFk8
uS8n2ZJKYUJxSX5Usvt3TYJMLV6zkdQHvltznYj+30S+ikifk9UuVqhJ82FKePVMgmd/xh2htM0h
xoDKxQt5Tf/dFVy3vptPp+fyWKNvR+N+vVTIFtBlU2xAQEM8kXkMuxCxzy42FlIIUEKJZUUdP+3Q
Zbmwovk/u6u6Q8zS8FhwUlOI89rdP31MApkrufbooMyVudOsxCg/t3UzgosFpmpsp+TT3ROhM2CW
wEsmDNZ8wkvCpncqraWAYig66ijTeGWaXLJNinsIMIKnDd3gxQmnriVEBp+MEE3g/0phDd98LxNY
RbvB7o/Bxv6k3VAdnx/pE4CJLB4ijBtbsxeon5LIs8Mho76MRxtOBOKrb/e+AtysQ1htPYhncD/Z
zkWHTfCvLiwgFMUUjQ14Z70uwekYyD9ytkeEeDH/ffSpzFG//9aThuMI80HwJGrBQNkrPrJT+1hB
QS2XjGXQSWRuZ+IoufVeIosm6HHMvWx6h/rcSLJg8tOr36sDp1nR8MzIKuzlKjdvO1l8QxLcJclv
lEWUJwQKZUCemDw7X94Lmxe5OpZwk1QCf4faqEF/rArCaN4wlzDkS5kMw+fp6nmI+xnNw1HxXGpH
44mwMZxp/3MuODB/kmmykiPR2tNxMjih15a65WRwGbsj1bRWms0F4JaJXlgkofzpRPDRSix2Cjlr
OIFBJaZuG/r9se3Txp4y4wNQ+eI4FP4JBxlYcGPxnz/38x1yfF194pgFQTEJSWnzZpT8luqDahhb
a3XqaqoBZ2/kDititLJwc1cEDkN/nPio9poafDU6gYlCPxupvS8JTZ/J4eqcShLmBazQSA7S9ejP
lswvGLwMwNMmfVs8mab2patoh+uDCoPN6d0CKoRWQ1GL12uNASqd7JsSM/BsOps8/P7k2OdLUrpz
XfpwGqVqos6DbPnVbfrlIlZGwcvkQS6BYhY/cyk2+c+B/S7svhBlC4/pLHBz+hpjEDcmDae3XBvr
ERUHXmmi197CetcF1GeN6nabu8Od3jgzt/z7WFwt6ncbA7+oYadhOVYZP03fANdbXHYrTpOx5Xkw
JUQ+Bth8N2kaPMcE0t3T5pzjlItw/Y7Fr4fp+uEnzRm6VGOCWTJQcia55zbjgTg5XdCGyy7KiRFv
1kghVy5qVDqc0J7aoyhzRlxjrNxyQIM1E1weBtGzoAZ0FkhURVnMadNDjJdxW2or/22WgAXn791L
1oN4h30m26MJjzARBtpWPcHeo4PKF5yEYpjNzy28XzMbPTeFHC7XCHDx2NfcSj60b954zjs7TAAu
JDNPAu2cwUAawFN/ZQoRfy1XXOwjbX8wg8qNI56tTHWn4R93LPADR2CHHSak8qIm7YKDQ/vDtCNr
DYHWKBLebNsJKqanuWSs6BcPmiCVNJc0IKNHxh9aNlWoKmYluumPllacnus8UhWNNKEH9qJ1jzb/
0L9P4PGyoA7SVNV5bfqAcpUAs1JY1m1cZVACKntDD49eHq1OCPLXeUo3JszXu9lFNdd2eUmW/Zcc
H2oWIyDcskrE0Tjsh7B5DXCUqdFcSuN52eLRZ9PcgsqeE+3AWd/mP3Qn853EnO/QmOj6cE8QqtEF
y8k52MHjtzuh/FMjkpN/RJb1IFEcca5/I7tDpo/rnKMeL14oN36t+rnit7jU7gLXUHuZjEFjtBIJ
WjA36s/9dDtME1lZ+DKR2WlTKjqFS4x3Uez94nc87E4ssVy3dHwCxTYNdxMoET4JQbXUOaPElsth
qwgBENNg+UnhLXzyKjawy1xPk1U5uZX0TQUjdwH0+nbHmmerqwrQpQyJiWVgCMDBKG68Lq/C4238
GN46xI4b092f3nkCw61jVEFoJ7S3/6Fli2mrT98aXmwBBau5XvckYdT/OhwxDXbZrLDIT3U4RxGw
VZwMK6r01TBPKpkqtfb2K3yVEve1VTusfMqOc3+Ju28qL9H2ovoNg6TWBXeIAFZXDUjuwrphrw1I
GYlGck4irWGnxw5J3R/vaAdlAjwIMg/+Aacog6GYlqnZN0uLxnGT7x5E3qi5dLGAD5GJuk9d03pf
BbCOZ9HEhxL/rxYHSGJYp39HhndrJ85zEoZ8ZqT2+qiqkjHbgPGEoPRStPlPVHt3kbHHXaVmDjxx
FVtpGd7kSwm1fxftwwuPYL9YqCJUgaEe1JYzdI6nXNpQtd9+yJWCRc1TBZYxcESc5saJAwuS+coH
n1Px/Mc15VXLuQOotCQCXzLXOJ0HVBoa/wsMz+7Pogq+iL7d4wxHoaH6DSipWKOvcm1sTIAovgf+
en0O3J+VwiQai2rO38UsuH0SX7cp8QfEGqzHLHOcHLQkOTbm5766Eh2Yod7CKTr21PDZY4gNlyS0
536JHdLSjFNNCcEjVLIkWeCmqCW/5taKbOxjF4F8Xr/SgGpEEIylm2/dvrdUt/nDQeqzrHD1KDe3
tIN3OnXEjdWjUeT3w3xgzdpEahwO2CcIk+GvhxGXhCK+uaRBpm18gzUPXp+F5jWOmNWTDTUOoMSH
c0/ZwEH/Sc8jya2wr10V4+1gzrUxuJ8+YEPBcBQ/qzqOnzkSEJZKVXK0VerK5RVwT5+4IMW0ni2E
WRLPplx6/FpM8VFTaE1BlDS6tD44yVOkTO2bTX5URngcfUw1BpKWzQCgTl8Vo93f4c35vqTXABTk
rqhabnMCKyl7Z6bl8lwpvLPpgHnOLhjg2LHRo4FMEHSmhnAZ0L5vbAT2nALzZEOz3LZ6LKidSWGe
q6rXFUCG0GwbnXrZw8mtwu6dOD5H8ll0XhCF+nbHRzh3vCqZvZRQpFx/xfKUtfvkThHdw18Oa0U5
chuSIjyQLDRuDsRXESmM1dgSO63CiB/6Dz4FYyXgBkyOEFOa6hu21L5c7gId7G55J0l+PbWpKqrz
73Ldacn9R+tx+CpAGm1kE42TP8JzDv9OrVJh+lxOztwKuzDbmfBG4WbGzpTG/6sDH3KALNgogBm8
rp++1//b1/64OqBri5+PwsJNwhNQTQv8zFUti4P8xobyvSF8f+FNJUWBIUbOqOKCQ7OX7ktFoHR4
5teu4OJraoB0Vi8rtQl+uRu5gndDXbgqU+1Vt+3eS8a4q48T4tWhImNc2DJZvAMwRtbITXXiwDhj
nvPh1eaVicWn5vX9r8e89uTz15Ap0ryXaCSDHaGmo4mqu6sdsj5dJQSZ/1eDGj40E6DE8GCk5crY
StsHayYG5NofhJtp4giwTaC+Fkvxb97TILFuCxe138wbGL1PvphNeVzfbLdhw6ZXA8CEgD3/rHZe
ooYBHRrbds6e+JtPqlKGggXNWryHfhkxdHk5RsjuFQJqE1hoMTYUiNkHC4UOsUcsCArqnbLztbVD
ePWwDCZrv1GtA8EInUsdvYCf12WePP57J0bP9AHyDMpyGemc5QBn6EE1TIK6O+27o1pkZYVRRcw0
Dec/1gsCQWaGnUrj2O2FtLFYAJtXTI35zNrOSrNlBMXBSoatDdaktfaPae7NwSdq8+rlXBnzXK04
+H6eTElklk5sVN3XSXu9iM4vaAwr+U+toaYaWCUd1NYDihnAz7BN6rZpmqM6pLDoXnmeQAM3UPZU
UWwYO5JrcRKsJ87CK11NtR68gNt38ICCZBfxx/MMUl5iS13CEqPubexj33g11CIGj+l45lwMkrg0
Qs8MiCFeq9fefwWSdZqKZrlWIGOoYYptFaCtvKZtL1yj/GAEXbibjpiflT7HmEO7bwnCX+0kz15n
BlI86rrernnEXnIHmHLNbae+vyK3T7AyidN8Oy6lZs5y0IEwmaVFXoPY3x1Wczna5GocnSEP7alh
f+s6q2rE9aFynjGCBb7Yf+94cdDoYt/UnTqni3IViZqZeTnIjvCd5PM5SLIAmwxPzUNe9k84BHzn
CqBHKezwazidD4wvF58xKJy+K5ezwLWdtg959TpotSEJGpbD5sud22/og/h0KSQg4BVwYAdJdNBs
gFp4bbupnDoYldnlJ7uVPK4anRhqzzuXZFF9uJZWx+h505ohykPIV6+Yas3nZ4YSLg+ag0kX3Spc
e3lm5xgJ4fziIAgEmlA/aXoXrvmYd3aP6TfrfMm68YEbBhp5//aOjAywcKGzhy+22ULznt/rHZUm
Em9Gm0XUZq6X8zNGsz2Oz8UzaOpYb1zP4thl0KPJjHtaB7/E+tEUrr5Fz6Fblf39cpz9ybfnJrgV
szq83vK5/G7hEsi4W5RWSlT28h0lRHvhwAp1e98EtxCDpZFWycvxPic2QfOshV03z/Hg0TaXePgL
Vh8gU5vlLhfChi5f7bu8T2wQuHaBQUDPB4mBcPak0+shsVHBvOHKa0+yZFRiloH2l+fczfVesuDb
1Y+dYh0kaQ2aq1hI2KAeg4B+W+Xj65xd/KAJf/oMv7C1+S++Zlf7mfzjYvLrpfKHfHSL5fi4IHVn
fBx8gWeVQnig/6n5fGuGYI1bHTrD/PkCfZwelx2+tio/SYSKVS1BlP5BM8kj3BXpcn6N+0qZ0Ob5
6bzHI4dYfY6AjQ3taPlyJLolkSG1ZNYM9r8+LNmQkIjGRgYP9P2dZLmIewH/EfYVBDjN8COCgniP
g2elv7nZl+DcE1bGVB5QNBhmGfFoZ5WoR69tTkxnG6VX/i86d8F1vkvw9fRV37URTWiVNDv158Pp
nE5QdXTfSyHkfdirGw9uSTzFHB0SeKOS6MveCUmCXeZF3lyaT6eukSYOngFgjPNlgRQim6sGC5uc
DsGX1K1PNADWCtidBXrt7yspborvoQBxD3gXy3+lcNR4FGUdID9pBYMzIKKUsoq//GmMT5bzUw62
2ttF+hZmePcGtz3yZWlVmHUGaFkm6D63FPNm4+1wXzfiEnWLjF5ANUvDy+WF6+o3Pw95oNbtJVW1
4MRQklWNgyqXXy8WCVpSa7hN0LemqHsPNw1yd3z5KM1mgvNugxp+sR8R3DxC6BACVRR0BDzbDkV8
6YbBeHNRTo8CNcetgmi5Zo7X5eEruoMpAJgXBM4rz5TFUMYNUmwxFIM9CexuxaVwfIFPE+5bYUHS
QVYkho6PzAae2yny+63lyQOBCPvbQfHThkLVMDxsXIe8mjKy04/uL5NCF689X6LwakzW+jslZuVT
HROZjumpCSs5b8bvT0zJStzlHrI41jp0VBft3EUAgXuvc3QQ3rrQ+ArxgmC0Fp0tKDWx9I2djYms
5piT2AzAtfEWow5BnA4cJzh5AP+4DNDmsbeQuW0PHd8eutH2g+ocestA6+OOsFOZG/8vGl1XD1DL
6G+FPZW5biT5w9lbGBCrkgw1NjB9BPM7NO+TbgJ/5FHGO5yfBP3LY35wCpHB4/IMFCm2yEs9g5Q9
JGAAx/JmUw0yhWY1+nfymuTwagCXmHeEbxRMeECFLCdtonOwsl+L5j6nyIHELsDVhSFMbb8VlpkF
MHgfzsYbPJ46c6hjJwis2zWiSgYQRPM3ATjWwFq4EsRtCpwLisyD7MsM/G0TVXs+2rcayehSIFb4
c3ACMUfMu/3iliiGIl9hpt+PckMPhEsrEnkQnNqDbc1EoSjygSeSMZTuDIWlx+cZbeelDWsKscza
F8LcQqettkBAkoTsuIDPBta7u2BphgsWqqJbpjkyzTzct4F4eUIBQNIxyi/M/Sje5YgCXRoUSZzt
mOrRMVswtNvd8s+tffxNd56FUL1JHR/LgnQXIEor8GjcnaAVMuwGfAofNqa6nTYfEZkGWMhk1asc
oVI+uzm6cHY8GMDO3s0tUW+6OQszwrPy2kirmouOif09WMDf7pMBKWCBaILznVV0tqx+VEpnN7iu
AHfgCXRmdVEITKAmiKlScaS+0JAJi1DIPOzGmYQ2mHZms5xFJ/5VB8tmGkmn23TUPCLe9sDouUru
rejHbrtEb894VSzQgw1mTwMbjgvGQgZtzQQ/6gRWM5B0dkR+Kx0JlplYWE0nW01ZWm5e7GrOtN5u
4xDkp1C7nn1Vbti7UDiUWu0cdzVSSD53MX96nB+AtzdaXj/+Jcpz8O3xWWgmm4EiRiArZL2bIi6T
lMXoLYH0E8EtpdIAiwu+PBIaF0hUqWhaP4pfRVe7rj/5uYg6CWw2tpyKZr4NGiROwxbpLPcm+x0S
G8/xsavF6Hwvr8OvXv55kPXr+bPs1hoeRCy7jzoE+XjsyF7Ez9JtOm6Oxc3+F/8uR5VYwLzt1Bkk
96B028L7QFm6ZRDs3I6nsFoh3PsOld/URq6CzjKuw8UWudZAf2USKiczE/t4sahGIMjZF4dHrw+4
GtQpD5Ax9yailmJ6B76Lqr5irxC9IIQb+fGbf3sUhhjTORjuVMKHooYAqcYyvOTZVeHUNkrPtb0v
MhdEq1diOy9HYx8h+cSQDWnltbS8dwvANQJGG69HK/MonlFx0SU8zITu7g0bdLmN7YGi6KkcILeV
5cRAffw421nYlPS7TeaADWbMlyiifQJ1DCO2eXXD/dmuawEZJFV/ItRuutDXCNgDTpn0/W52ndgh
3QinYuqpxNWrMdqU3xVEvOgU3CTFQYoOtLUKBO1g30A7OkafY/wGJUGmHW0ab3Noo480p4UyswXF
z5t4fTz//uS/RzQhvj12z3tC4aIcNB2d8s84AtJuW2PYiRreO8J0jJDtcNJ4ECFrP8eaQaY5U3Su
QiWJIAxeI/3MohkurL6WbWybOhOETn36+vrINMKPhjB6AffHEIaZwrXM7Gyz2iXz1UJVnVMfMDR+
GWHEtncqUFiEWrkzJvFt+vEfCbBq3fwHWMbBnRTXBbImmz0GB4ZfFXTxcHk1uq+R0ApV0Y53o4qK
3+YVTebpXS42n+X6A5RbK02Rnngg2nwwEWqOmd9ht6oAcs3zc9t5MXcSHHfDAl0ZuHqIHajDmZ4+
FUTxWm+Cg/uTFI/EW+Ry0arTn0NRPBl9re4LVZeTTW8mS9qsnb1xyBvlvq5nak4OXCzcFliIu2Bz
pO1/yBsG5zzd6ZNSfg40LIE8j27fYiTSrRJbEhLHsfCSM3RFUcS7STAsWnlbcl/+BcBZ6OFRFADH
p6J5UTwBVELkgTLWpd8CiBd8YSiAovMQ0lNLjNdw5j2V0gfoG2D6wZhMO3j8gg8XsJMnBwx+6xI5
huV/Kol3bzspL4rtlhsUkoqeSAfojsAUJkMkk001Ip2fMp6jOMGBAS9eJhUnh8ZMK12rqtTg4nYe
qMdNq5MfF1a1SlYcUuFEp33TxQICyjZzo7hEH59wlIY9kOBEEoxKKB3Mh1HLXTxnuq/seDsHOeTw
VN2G8KlJkgsb8fb8FBpSNuaDy9d5JcvrV9HKzTic2ofJ7zN/QxLfF5AX0COmcXev3H+Z3zBK7A1D
3ddt06UEZGOgdO+Dd6jfHpuPuNTqeFhyppmcTM3FVsoSOz726KeyVaHeQrKwiGQ/a+Onh+QGuKri
EtpSZIlXnTeilBmT8SHzBk4MA2itnz2ehEJC6t0bmJAtu4O2tEz8ROXrM34Hhl/irI/o/ANdE9Xr
e+Oa1ri6YVv5mrrhAg8DP5d9bIOs3WozJPwBBgIqEtX3jOTH3ODLfDSPbvT8IA+pjMAeoRrSnLTP
t0GCDnLHepR02vHczG3tibUWxbMbVyE3+6bnjYpwmFt5FZUqweItZb28D7VLjI5+oOKXEUiYRenq
jFXbSXb4RsamKdouC/zES9sPMwC1yLnwC/koJ4+ePAEeZPldi3JmBMyAPXTYupgMbCwR+33bvAJi
yMEdgaadTPfLjX3gwcmmaWTcO3jQ1nRMzjyNs3eYE4ulOqTFCAanxwEySxi6lsDsCrHVUwoPN/R1
zD8V6cJO6BdKwGHxJ2BCWlvzsjBMvUKHKb0IsET3y0a/8jEhXXIOyiUT69MJ2M+O8mIUG5ndqZcp
J0yoy4DN/YNMZKekoKsbU1VBgE7BRGKOPnlTLDteJNEsWzq3+rgkWz9oJ23jiR67hQeRD3b/xkmT
DTm/nI2d3ivI776a0MZDvKWX8d9+WUAjF8VmMdv1WD9R1TX0m3XI5yOvnjnw9Qj85UhX4mUcQBge
6sEq9P48eBvtRXsqPPAUL26I9D5TUWd63TQt7UkNtJS8gB7URYF29wLkzs0smd68vorurI9R+zYJ
lZwKwNnUUg1t5lD/WzuWc0Gmq5KXO1qdDkCwCz/HR9nK7O+4rVnjXE5IMAeywF6JKJI95IcRaK7O
z2xZRQi6hmZmEh9q5cF4KseyeWkznTeifHj392mzn/F9tABeyeKVklZmSgAS6asqHXIGYosItkKr
wfs8bCKY+yh10v2T9JEM/Jsczi4ojk+5+/v/f95EOzXh2M8soKhp0+IBvwBJGCshYRNLJ7zRPL7n
Sbp50rL25VvCmpbDOSpCRX+W2eb3LIkN6OOtVqvclrgY7Z6Uasks+h5Fl8blaxjeWEyyiEjJ9VDJ
FQfXGk4RidKreTIYEy3oKsRasRsfuQtV3gXtuWM7FIbjPjzG4vjTL4OSaZwgc0gDW0XBqIofaIIk
iQxRQMY2R2ZIvtj8RYjDI8LEbR2e4gBm9aG7/o6+eNF1VY6gIY6RF73mQ9Wzbsm0+qzecgUAGrhu
RMovV1KRptYxr2dtpBpWTSZCW081Hk+0ow8rsJvOn/cYIiK8GAvRTIRZrdKWWJzmhOVyf76oq3g1
VrbWmghbu5Lo7i6/x+fKw/y2PDWpExUMUjUPGoZ7owxgUPQixbcwJ1vdpJu8zDHRkUVaShA0QScl
C5+Ox9FHoCM/eqe11rFXa8e06wTsG3ioExi8p6L/8S6VtbAGylI2YEkgz1cSDXzNDGCMcWnHdyQe
O4G59LHyz4pv6kfF0KEh3mCIHOQIP6b1cC7ChBgoYBz/iI22UsafGSwHNl83wNBkkL7L082Mc3Jg
dC71bWqvsYpH8ZTqJPdaYso2g1m2W3IMi/GRWlcCEgCHn+VhfPglfx+E0ALfuuIFfue0RoywzGJC
Brfw7i4OTJzk7DVXmVkaDqsCjOvUNSncedy9aBBSkPOtqKLVbSlz8ODmgZcKBML+lQlnbAhyRjYr
k/oe+5xwW2YSAvwh6/z2NJueF8TWe7HxOyk5dcTwTArXcW+bUKMv+twYKFE8h1ya5VeEG8aY4gt9
yTWTHZmTFJIyxziyea7B25kclRst4M+Ub1XAltB2i4gmi6NsMFFCLYkmYFjTlbIErVHjQBpGbq6T
FdBxnf8ONQ4dZrkWERx/KWbr/C0Kyh/uVFo0fMTu0vEGIIgJDy5BtFsVmmeNU9twRS4nTMjj/V90
ibBlIOpaxMkGYx2QnYd7meEg0aqKJ3nh/QCsmc/LiCsoxxdO8iAfN0cDRW6F9L8v1zBKdxJGkIsu
7Mmjk0T+uMdvs19KnzBVS3owjrUojhpsIb3snMEsJvxbF7t5/W1ABTS7PjKArklBigHZ47t987A1
vv6MPtzBqyUX3jqDS6J8MoSDzKn6ijT9pektFPYRCfPxFXcWC7FKx9bIc6uFQaJ7z9f/ZZfENWq6
uJ6SqA4+25AanJXY8CzVeNoPngMb8+sxt/CxnTAErprcfpiD/7mRkWbiAu2o9RUoGStGPcTyok71
MyAbiYwI7/r6vwHQ5akyw+NEy5RMHKKdVhP7z9EnrPnhSFZLQ7zJuFzSprW0LqaTfgJpSnxy5AfW
6P9vAIlZmFmt0FUY4zWWNTKiSbeL2Et7NKl4kMLhzPZrvEQd+uXoZZ/upGTDqJBw8MIDheb0AItW
k8pg56EX5i9mTJtuZvRz/l9inZ9SmPTQaXeRjJo7XYaRupJriIm5dLqTfddz2wnMP2TlkOCjDuHz
CwrE6gUt6kAbH5FZLuHVCYKLgwQWEupTM55wHtlWzIDak+XIGYwiBIiLxRpJ3vCEhsuGVEXvrJd6
LumI3BXYX5rIN5XJ4UEEKsvswFKMWZcYUib+wMGbP1xPeHPUCZf9kwMVl5V1xjE+PmSD/yF444Yw
lIbbnXt46VX0sDuh8DJIQzzBN0Nxh8gF6pQgBHwxVIqQF6PWTspmWMV0FxImjpZWPtTIMAL2h7U0
FmE5KirqXYPdWdwE5c2NFlogpU4+Vh+tcGro38bOY/DvP4gTuUHjovyehAekXe02T+nvTsDEyvFP
PmJtH7a7JBCFOPjFn788Z/IPsSTEtkMBdW7TcsIDARWcvAg0Xa6pw1BXy+X4CrdHM2hckpmy+xY7
tD4m7PjLCdx+zrgMCCVVFdIqL7SmCnEIjFJXAXr9vrpAtgOkPDBFhmMR4zFoCVWExDIa/49Mqp9p
69epmnVFAzmZPq+5ocbtYzv2REqSP79bAul/nQMK2xZrT5F5eCMtiJTdFm0NmDjifvmRojlPnCAb
ImzIAhd80AbOEpTEba3xH7JLiqjxDqT0JfOWY/ViyXpmPNiE6a2opNaE6J0WBrli7g2/0M8OMDar
xZPQtrKzT5Tr6aBFCiNR4kC9Rp3A5QzwzJRvKvtd/VvzpfYbH61GDybKxeAy8kss/KS1mlPETFaJ
hPWKjAo6ZsQx4T/J6ou9KQUQ968MY7mNZZhQQH30suB3nZtDzK1kKRthQhj91rjUQ7Lek1WdJWx5
CsZho+MzFFTSuxMN7QRspOPGbVXtayk3POD2gUXghweDRYATYQ+fY5JSF8OTAsW8BFFmGAF3aMjE
28ZGyNEEoNlt+e+PWykFsF4SLjlHUIVIAJqiFk9N99wsWzu+CqlRlVsQqFLJuAc9SdAU15UDebFn
bFQGSA+HDL7oAkWhJsxF1IN9orcf/Z4KBMWYFQmFFbcyZ7T8MZKnhv7vs3p9vdSRfJC4Z+8Cu+TZ
u4r4q6/C5WSnrdwpkmAY2Op0emjYqDBQf+S40hN0G+1Yawj7srNZyS9vJPxJ2RMu6NSA2lO/M0Tk
8ZEOrk8xUJQuSO40/dd1Uy6zXFLeQUA0H7qFqGF8UGVX/2PnicqmgpCnCBUx7vHEpn3R4dmtjOb2
S+AR6fVX9OXIgyx3UJyg9ysmUlTfAslVZfiDKiT8UYraFZeFYcJAccLETWN7SULdzYU3o2hSdPHN
1osf5EaIXjj8VP/n3mBvtnq4HpAwODHhd2ThxWXp0ucXlStb9nS8rSr4Y4ukcwO1k6ff7Rs/YTLd
jfoi4/fhGL6k80qIvQyWsEDx0Wao5f6zqo2HDxLdjCySFpBb+Hjp0U2Ogw56YXymaS+mOBq0rFx+
UDbcOMOCCEvXwLF6WouC+qJ90Pgrbq/0q3p1kwtuEfruJlOrc+gLn098JFlViIA1EYfh2/ACImX5
68og9K8c6+7hf0RIMuml+r5SSElvVJPVF98NoKFXxxpANjNj5jWwMXnv4ONoosRf4hB436BrdW4e
JxG1bR26Uk9LqZRdWYpEa0zDobMAxSfTxtWVsm5xs30gi4cU+JVN0k57DpEjwbGzVZrySoaJ6qJX
viVkFQHYpMBHdr7N29TTm2hHUzYL9EXp9eeKzrtc5Sb+5LktHrNEobTNNEtJdzLTIh1oCUaD+xZ0
Z8Jdl+UZzNa6qlTxIoblRSt6N2e4JQEz+uhmUBU3NKf+6tstSp0X/mHZLqf6tJ9U4sA/U+Q4fNmy
64tQy0CiGRhxw27Ioa1h57zgULb33x6+wBSHEqGYYD6jY0iQyIoe5DIdqch15hNAbjP33xC1rdPG
ytl53V3d+Iqh/7GOfv7+2LLdHMFs4b5Aum+VEiw5UM8n4LV6q5mZfJXHkiVHh2/zFNVSPl1UxzaM
DTTJdEEHNTW/WzreXxEWdTHkT76x66rBld1BBhqwp/aydekHVXdjLdRnRnSglbfUatc00QtKSk0f
MCoQ+fxGLj8OzUnKvCFB2qwvTlXkeII4abceUFb6Ac3nXePgs1sXAmBU1fLlpLLuuHo5fpr0OEuM
+UUKaa3R3iMQfNTqcDyPKy1VP9fAUsin5C08uSPc/5JmFOem1tkOFF2CEFb+FNpgi/kxnmc6RkHX
iIZbLTxhlHgJEbl63nWgdIlpTLeSzYjipHXT3wH+pDU1Wffs1lIYGZbkS4f9YbcXVHmlEuiEzzQi
liwyYyd67E/2oBcz6Ugcz+KdGP/8N05M55Yjo9PlP/PS9okOcHpIpboT5a5MF1VKiSMZ63mT5q/e
kaOiXweLIgnzSbEf9uyqbhKDEjTudaBBv0jKtb3Xn0oiJ0LVtzzETF0UO62n2Efza1h0NJHISv+e
SOiKCwI9YwriFPEIKa8mqOrfnVqQMWy/ixNakU+WrORN1qThI6tH//EkrI8Tp11b9FAys59tK0TV
O2TYFRPn5cF2xBc9Y0dQ76+sH87aRsmKRhq9GgleHtTLN7F+oYBn8lcdsXqAtfb3RqtJdW3SSKRM
WGizuH+hB4+MnAgAHxGRJNDKjeoqGNkbof7IvDdHZw+ZzCllR6tHnPdRmNLQqv3th1y2bQqGRJHp
DFhsa7aM3USeL0ZWgMsOpBP1W8+xcmZnP/VJRoXuF89pDFXR5bINZuQ0vUfFKzK4dC2mU+087pHU
B/sQpeYWptzt+5Vgd5wE6l9eEbbDtrxKOHv24ON8FnxNa4hyVgGDZu7i/qC1JwR9KURv4QjzQ4QE
uNRH9zZbDs1MmQWi774LZrEFcXsb1l/1qWfS+dWnweFmOFFz9RRQrDNu8nwo/LZN5rkWjqUcxCmT
KDBAzMtow65JHoUUH2zKgdpfn1eAsvlQLWiMnfU1D6WWIeWFqFCyehHumRw3nGcBZxQs7p8SVeLL
bYQMsaqs9DEn7aqFKfduyKB21CBv2IuxcH6q22g9BBeMvDsWW814aIj8jGy38Bb9HwO+gyBUodWN
LSYyYzAoWgbC20Lx6x5xwtSVh3AgN3dGn+WqglWcXd9mdGzXb1e3ZLePzvWvn5mhoA+UXnmmxTxN
fN/UmReED35dyxyTua+oBeU2ED5GVxTMDsZHYO8DTfrloXweMOlP0VCPFnWiUb0rwbjaZOZalqtB
9n2l1Zi0KTb21W1OVpNZdMTreaKgV9GfPQ5vByyhV2Ew9if6mXpiNll58wMr65J8KYODjHIc1iCh
wj+m3dyfJbT9+wPJOR6Swj8rstUaB1NURF3BCwbZKxoi2VVhYO3vJq298MSjxepCtkpMFRspTM2E
zrES2bQtr1FvgxbiMWoSWj43cdbcaq5+cZeJYk3wcO8UDLLGJLnjFJ3I4cdBpV6+WWXmlRwvg7VS
lOEoJffelNHZoUTj9Psk5qSlMPeaYLazi/iZaSiAij3hVTVyhWeQ3BBB/YFOVMArHzIlLpQwGTtn
TegYgxdrMBKdNNb0rl/j8zfLct+s2ITg6ppzLziQe/JyNq4QlW7M9yUax3Vu2yAe5PSFdnzz7QPS
qD+Uw+exXy9DX9CvdSLvZhv7xkj0HruN+G+2D7tU+bwYL9q9U+W60dUbXsx8RB4x1b4mmwwgIc8v
KRx+HL8UKflA1aXjRWIiGNPSuMkom/7UIufOqVHC1if5f1E/K5ZB4RXf/w5KIQlsywPWzXSVexPy
hCo+KbHeqxqyforso2jA1TWMtaCUZCp33ViR0VnxjLDWiwRJHVTgP342tOlUwFinQdxM6JL8VC0C
xCeoc2XvioAJ+i/+u3t/Rsdtp80bR88j2FwEX6Ju6/w/P2istqbB8x3N3oiJwqXYMXF8QySoAneZ
Y2LQQaHq/w87GVDJLVvhjDpmUUOptbnx57w934ul7HUNfLatca4qy26nk3GiA65gJ/7aD/JN2vMR
WbK53bVFKu8hxk6wM7vVNSyBoBFu0//Gmyb1VV1x5bjF6VTh89AFsFqd2u/Nfs4iwvZNduHjKpri
EgevTf0aed1BhoXZbrHMst4T/Pf7Y6476WGPHxaaCclILXSM5kBaFueP2Y1SjcOM17yDKLleJbjz
pH4fBH8Q2U9qsbhtBek9nlzR9+AgFndqBKrGJ3pUG7fQf+rWYfrPHQVtl7DtyZYFI2Q8bL0Hmxqe
hG8AB45U1fwJbCnTRuGD+XXIUKcgcVToGal2Q/c/er9W72BYb7xriwgBW5CGRZt6B72VM5X4d+WP
pEjuW2zl0if+tsT12ZThqedPzKezKVgT2iVc42qWEEgBQFUKhaxKj2dAv92VanY3JGs3mIvmOY8W
B+M9217Lnc7j2Ji4brl0vVKyuMzwxP8CaCK49sP1CRTBCQnIM5OMBdb/BHRpjv4w6w8OEp57Tljp
4NHSB7R1x0rb6L7sJ4QsuDs1okMzQ0XgEocTsgURqxGGAAz4uR2xNClQnZIiPnrxCWszjuNYHnOU
l0vjf32wABFVDU56WNoUNmtbbkgEsi6EaTgzhLTCENj16Z2y5kZXbr0vPo4+GH41RnghOboYykVk
7+w8jST0r8H1w5jC8qVDWCfgO5B7DdhSUsRIT0NnadBPB8iWJxMiGxbmMIs1e2vqGWUwaV6Dhy11
OIomTvUL0TPCF+z0Dxw98HwN2hleBPJsjRdaT5dQHC1d+6KiggmWFqYRvsFYa+6OWMuT7FnOMCXZ
DlZk04PGsThD9cYhPxF/5eyPFdVe5v9IgsouFCP928s/GgTvnna+YlrtNoWjAktH77c15OMUun6f
D24LpgE06bB2hdi252/XDkivWiZh4X7RcIs0m+y9vtEQhxxbAHDClbjmQB1s+GGSp0K6jfsfbL3L
CWZmVXgJ9NSqg+Dh+NmLfqF2MjqrUjip4HLcfkhlqcFx+d5sSBW0c/ML7Sr3ljCyvquV6VoK6Yyh
ODewe3n1L2ap6RJHNg1ta3Exhku1vyq/hsdmYLmg9T8IpKRCR7yYb/NhmKtcvPMUKJfVsqKTXiSc
dvTaYSV6kt1dJEmogk/cGERwTJKTyFywCdCIzR0zRYrsPO5UA9hkhp+s4TlQ37Cc1qyY3S+BQ0hC
702tzIy7n8JoJSiC95Tt6/7AUKquPdAhfOijM4x70JsSJavDokXtuQE4phYpnexJlGnSehndixzc
vLA7Lp4gHHps2YRkf+WgAoqjfvQKmSd2wwZBK6P8gr3NSowycI7boXsQgd29aQCiTmhpMF++Nodt
kFZv5zHgoagz3Nx5SyGdtKSkYuPKfdIhgfhYVhXNVZmEt/8l7cL/mPshItrO506d32bZIXAFWmdn
4LDifUCIdOysRuLL4qA4eKU/5vB42NNJ38+7oczPEuKbTNoYtAMVww1B8cM3d2ljdDEkVNWOkkfn
pqxDUvgfcFiKcuPqNXMKPJtVXJ1bzjeUtUk3lG5a7nhRVXNH8XcTqcX++htoLMoXYUoPMOVETurB
bhDT/Q2W44LBeuglku33gIs9PcytS7NW8f8131NefcYje7w9qNDQ+pJ4eQ3lMG+rt6xu8HyrW0zZ
eI+1xKKBAtDqlLm8NFe53RwxaYGSDS5oKwuw7p5XOMRrNWln/wxKfe7bMwBENNy6zx7YREWfMukG
LZWvUcoIm+1Ge+gGBdx7dtMwgWM7Qfu0CR8YdUVpoTwfVj1KoMio9PUg8Xz62A98qj6pgHRyzUrL
tuvTLI5e8JEGPdo0v0QeXuJpzbrUHcArYjpexMhO8UnAk89pWShWdhpfr9NAuLq3nAtmCjYYCrba
Cv9Qbt2ZsgpV623GNDUgD+ODbiT2XUsjOxiBsXZrH7wcLn3Sy6VKS9ZYu7Vf9A9U+WECcZZXhYju
QkOn0ZVZEBOKuklciUc72MZxxCI3cB1id+0ipOQorhNilGdOtLJMTb+YHQagXgIhq8DW/bMH0yuF
Lk5tvOd5s6Wk7SIBT3zWMGbLj/0q4zD28I5saP0ZvB+zHQTwohNIv6quEig94bpiGApaWgQm1gao
VeocWbQMBHRfFz0Lo4IZ36lWAqpBRY3dGqWDm7HNdi+1dT7ort6wen/6IL0hjnvIEdImY3yPsiZc
u5WzL6EDdSxicL9VllZHiK9Jbr3njg/VumjVknbEslvV3ha05zyaHnxBdlQVACtK1vefWE5Fr34N
eSv+FaHWJfi9C3CBdgdZdjL82odj/OgNfpbFodVHBUPByF2r3wmNOoHyLYJ2zmwnEmVPIKBzu7Ho
HiVYRFVbRHoEpBk3vuGwjzwlA2i/qzZi9kUT7rraC2NlETU8dX8E722z21cs5yzGignTkLBAWeTA
0Luv8fUNbnPN4UdRjstk33Ulk6IFbcbhLf+QUhoWLQUL+pOZd64Zd6IUqu0gUu9qm9MCg4M7WNKY
2Ife113L0C181eqqKPjd2uHkIrh3rUXQzYM3t8LuQiikTI7CbIWDDKvkgMR+AuqSC9cu1Xl6cUHh
Ev6r7P1Z+aodk+RRj/l9T+7aR7SzNU0To0lY+lp+PDvUnBbUvROlXDDKOV97oSvVoRRBKf1fxCL0
PwYdYNTiKchr9txdFmF4fmHg4bZmFlXnwEh223yIOG/LGNn55rt14eAcv+B8YdhqjNmbpgHsIQg1
ehpZRUSs5NI3w6LfPdCNNBF0mjLRxYFdyMiOeckxWqoOcq4AXWGaL+9Vw+j6wn9HYIr60dvvDBVB
myw4vua6bnacYOOFktjfd2aoaJRc8Ulv5+C1W9Qos9DIPCb9nz1rLpHJ8p+QAzNMqizKDvW9OKxe
Qfq/dPJGMUaeDr1mC6N6QPEzOUZ8J43UJv6OU0yrmdRPuYioLNxzfUCIV2xW6TivxQikI/EKk0EA
ax0CNx3mV/eU7bCWDU8YlyySEZEf593aAk5dZL6YmjDymte7Ay0jHFNWtSdCSndDbVsZyD5qA4XZ
9phmBLGUh5zPw61JZuZ1c1PyBZBQsV/uuEsfxsWHD2Qr5cKhS8+UqKy3bNUmzTHxAhVhuHjB/Vhw
NktXQZejZVw0SAlDRkJKJ+ba5KC7+QYW7wFNuvQvVRs7fe+XPTAmHFNT5/LqpyCin48lsPR3HqK6
vp81jFssIWqvtjpNsrWrI8bUGykdyHUK9fdsTdjWeQ1Pw3KlHsLwzbyaesapgRWPXFG7FpFCS9AT
rxovePlhnmzHz76ZsjLUfCMeDr3tT7AOrgplwm+bC2xXCdHofkif3/K1rXGgGwHEAEG2Z55rvvIY
8qQ8HhGr2M9aS/YOpXfyCViMS/2/AQ6srdX8TMmtrhDg2HDpHvy/RqHJwVL7+jXb2wZ08oJb2LCg
fF1xqrcR0cNkChqQmhLqfQJpt/hKd1v948bgqOIwLVUNKVB7K6hihxGoKyvtHEhBy0faZDHuw5Th
UbUcIpGURiqj3qorBDYEOM7UN7vQs89d3LInopLP1wEJZndSHAkmYEvgKzYQYulS6MUysissBWif
eznzGZVDC+Mb6JT95XIP1Mf5BHvfdP6cGoz1SJjEe4QWbMo6nB0zeRBpnXry5p/ZYOB38S3XW/QK
cFcniNfU4GgP0ElxgKeYdSClIjgkbj41+erWy9F2gnzivBfTeL3jDVco96iZBXP9Uui7ZsKdbi2A
Q/amC7ACfTfcP2DY0janf6D/FsO1GL6B6eD05mR6Wb7iX4RxsSi83hUmJEu53FQ3OGFhoE+UeAWP
GDdIUGLKkR8HVzb2J5v4VWGybTnDTYbMQedyyuSPsLFEPfD/hCdNoZsZmUzIM9WmQm7vAIMk2fuQ
E/pLDehOknBKBThRKtnfU/RWBeUsR2iGrsjSV1pgR5JtEFxBJXH/PJvvECauMMHDvo3N3glyVcHx
K4cKqy0nu8r7DTslMZgj570Vjagj78Xza0YB94wy9t0mkcfO7kt+Twir71xc5+x36I7/TpvNKNhp
4ZyZ22gC4cGjFAOI1u8KWqXNpYjbQluDKyVEETi+SsuIIc9QncMLAI8ttfW5IfILWKPYoKuloauH
Ko5uHyspKbQhxsHYrYy7LjVeMQ87I6FFcJmqohfVXOxGKWhxPE3Knna08l6CmdXXtm65gZfP3CPT
nFrZLiRiBZPtiTiPSz3FaMKEcbG4yGs4HI6oWcjTKb0iHjpnbkIxFqlKnErBxLNmr8yiqPrA59Jg
rtUTgIzhN0o1hBJM4xh/YjcA9cwElBFnfr5TZ1tAwT/yFHTgJHF2r5Tda2KOgi3ewDE0bL0lxP4S
k2rQKcG36lsWuwGskU5PI4YJEgaC97+cHeWnZ7uDtJlKFA9UcGZjrLDXRCY1rviVcOLCJlrgvUNF
JuaQzRjiU0YJynQS7g1S5EW/Vyr0AdlBrxstLUb9+Q42nhDutG8e9ZqUmKwTn+SNvMb9wFKTu0SP
r5Ps4ygp0w9kUshJDzHwcxYSvhk7JExGMM7Q23yK3S5ZVW/XL08nK+LPjsDhuoEpg22ISXba+Z10
NzaT6asxhhaHPtspfHmAmT3HLsJ4bNNrgfEFshOiELdr7st4euqYsOZt/bknTGpxOSpbJQs5zE2M
Q5oOTEuOWLMWvTp/HuH6NDu5vXDJPSIH+BUT01gqWUE4YIfNN9KNB0WugHWjjkjYjhdn6tto7jX9
yupOgSvA6jpN1MilpRSYcIOaL+La1HaW4QBqyKhmrysL6U9VRQUBkFD0An45FlS7QykCkIwshGhE
TXTTyFrPnDeu7DdN3WJtIf8Fsk3smRoTFnPxaHFZzm3o975+wAaEHrAvtq98mHjMJv2z9TJi8/Ns
IsQRjZFNQZBmjkuP3kmGxmscT+HntRtVmKqOZeJzi/4P+dzjmBFXthY83czzoCu3iEztmu9MNQXL
CljKY0AfrMybhwJeKorloAOkQLZG4GukNg6zYnH/zYliJxfgFNjPgbc8SjulHTKlYAtxdayH/uMk
EPkSeiBK8NFTI6aURM7ptz7xz+RYJohVyIxsoRLOyPTAoAkwTQF33ixn38+h1UFpr2kShwNDjCpv
0Cq4/niyqJlKM3/UqCVChfqgYVJUpjrK1/8JkGmAn8rhEvNtBfW9vlundkthXOLHvYvr8sC/Emy8
dJiqXw5ZEEjP4PZ76E5XVZrZGVe2Ot00up+Ke7erwwfAyLlXfXfRVb/ntkctiDH0tadudkJTE8Sw
nHZ71ZzVk/yoTjWQc/TWPNsn7QJgBmsQ1ysTBJhd00OJmN1pEf5ymLgyAWD4R5mFGxJA8Ov/L3Yu
t0GOvByBYiiLumSAwgfGHYCNS7dq9z9rEtCeJOEUbh3iX8hJztVJ2uH4uJJmDha/SEqKBhkS0Xy9
qigxGIox77P0au6SLmwTQblwuMqQ6vQe9qqf8zOwu9qj/HjvPuWZnTk5InFsbuu4Jd9CYti3yW9c
ASCZdqEVrNSAA6D7+PjtxtZQsePJtS+D8BAwHgmg1OB8Wp4IC5b2dobcS0N3dmdlX6023Uy9v2XY
G3zC5mQa9CnjsDj34VqBABOEan25WHsJFJr1iO71bUuPzo7XUsvtIAkq86KpppRMBaAGC2NbvT06
V7FwYYnsM6EDSV2nl7vwh5YTAS/7r+i3Ka0LneuX68ha9k+6AOD94jBamxeB/tjQ3Hr5apQaCIUO
euLq1SZycOufTA9yRko0wV0XSFCT5d0bU23Cfxdw87yKlXuvRu5a/rm6dR9RauKkpXIa7dFpAJ3r
gDODZy/vyT0hHNGU9IdTHy/QkBEf5Nul2I/iH528jkvmyoBxWe73uw71uoK3uQ7f0fmhRMHAxxNg
0S5Sd2dMMOzBOOiA8AM/BMr73NqvC1CgG5zVNLydN+6J7m/Y8ny8KLbGMhH369c+BHeCzmZaZbLZ
T3bhnXRf4U9s1RwNJ/pMSGOZ4PTi15Ha9irvQmkfvEp57lqXLuiuNFFmMtLuZ54ijbwFp57tuz6Z
Tieb/ycGLvyemGAjffZpJT0eNRYf3PKESDeAuO6o8U8Kh4TjqEbSOnmfmrWywAwoa2ob+D/+p3bY
5GmylVQCaYfcoDO1F+7y1Q2Sg+g83NVezCjTDecGZ0uY6nYif/Auu1z/tMtqozzqZEJmc5oLwIVH
cVW/zIz8fi/40QCA2mQydP8WEyGipCDuX6Dq6u7oXaEjzZWnD4PcOW9EJLo4qRKG/fLhL2+liy/i
2+lMjFGqNPBJZJx/caefuk9cfMqmgfgtKa9EmAqrSIff93IjEwbK5+NKO5T87KEamzLyB5exgUop
fcyzWVoMbQUST47S6f8bv8rzj2vBgp9g0GTQmcYME3sEVtUS/AgNC1ZcfUlqS8L34nJ+FQ4gY6nO
JAMHir/ZaiLkGWulbzGFv/5rm6LjbfRfCMm9ein2z81viZILH2sKA1lV4OUyoMBO3nQdwQM8+wIh
Xby4Cl9HD+FcYsszFbQkLK1eMhxoyQkQ73Hn34Qj3UVHyQdBvfetSqXqwFrP69tN0hKROh5GN+cb
z/G0GI33fAtwGYFME/RhhcQdc+8gzg1oXCapdTQUgJRhN0YZrGgVRBr0wBamlH5r3U1MlYcDO+kC
JccEXz15ZM8RkQ7VPirONquBKGzsvtqn8qcfJU5j3WsGN82KF3JM6YfZxyugqeg6/a1apw0wIdGg
lF/t1xySwfdYLKsyP+TOg/wdNy8vs+wame4WZKqxg4363T0cNvzmrmEoMra9JW01q7lKJMZElRfX
eE/9Q0mouqMFZHMR0sjtTirWp6FXbEJFfTv0ENVDRDSeRwZqM62H2OIDpEt0GvjsfTTiQeTLOT2W
28VjUbwmwTpF+XPh65y3gKebLcnRASMTaqLzMo+rjjInFqm0N79YGSZjxM/4BulG47pQYwb8mNKP
plKBe2D5u/DffDgjyCoRoVrJPDuQsVEnj4ygtYJh4p2NwQy4yiS9AbukO91Nd/u0Dzpe8RepO9HQ
Wv3oc6gXAYSDEgqz9O0sMswJjna8iWGSjeJwA/my2eKgXWaGauNmAq9zM6DAZhdb3zV0TnDn3adZ
1urYo/Pvn2FrYqFs//4Xf7L7ZNtDwctiSe2W6Wd6joytAtZMZ9EbTgrQQiZ2yWyt4b6AcQr2EMfc
RdZH9ndU3H6l+LB63RW8dubQw5dGwjyD4bfkuYau+4GMxa9dKFdjWApJBlzq+ppCy5Xz1n8H1e3b
S44SxaaQgt3sm6dxPhMJN/vP5Z2sr+HTW/nhES0zPpVJFNwui2KPvjIbRSSHEWT09T2997lDOxXG
fHwQ3RT2shjCFzas21VXS6aUtlOcRFQyrLVzlTKx/ahsy+QaWuOePHhFeazMNz/hX61h4KzjYxGH
RrnYJazdmGTbu+fJvrJps6RkRCShf3BLBEL+mjqyeCoVH3LMfj0SEslvDyTal2lQ6qNDF7ceUcei
6He+64IXzy/bUZnpNUTuzOyrncJ/JGsfvaSdvpVU1hOegNZ1gly0YHJUUMPHDuP0eJuvauBdxgXH
RaOsnIw3uEwGLBLxrGoi/sdMGb7r0f/4nGBOpuVLBVGNsnLxu6OEyN7mn2tzhCgf0VghMU/E42ur
oATC3xMoEPa0VF5MBFBVZXEzdy8GPIoiOUDSP5mcX6sY+UWACd4MJh6yOpdALOFC2bgyk8i+23tt
avzG5xOilct+GRGzfEX/UclEelPTtekBow2JKlJzSWUn4RLcZSegQvhL/p/QDoBuqXzJJ343YDaR
MjTVa2Q2deFzhrB+Z73xDFxQs9++3M2gqBwLzJ5FY/jd2jQq3JI5jKQO7yHryrsljVomln/7TuQX
JZByzQ4bn/psTSW0sE2zmCuuhirkHbrUbXA4T7xIbTANXm2BcqHo9Pu8xH+CoMLnLIv9CjqXiSlu
4JqOvElgKOCj2SCRP+zJiZdrSWNYxj4Mhx8KLYf2lNZvUUrBmyRMfKNBhFdQ+HoE7kGtCKcq3Kiy
NdEyIszsmXzumZgkFHvXQoa6rE4r+78rrOTFh8UjCF8+m1joCG0ax8pUeY50ZSSNrkPBnqcAtayL
iAVf8RrpgWG6GhcoamIC66vCs6NPbE1SmFrNgZkuIHpUpR9WuSAJ8IET2ClBD+vU3BPTgW0QKGsJ
PmDEp0jr9LwBZ5p8E6GjkmU6Yg4WEtfSzyiGGqLo01TYnDPIZwyW/ndsc8INIkNlrSzJb8tjxmBh
zoP9Ef6jjm1MEjoqMsFQ4YTP5pz0oRrgUY7nxS/sTOSsRK6fzNZTY6wEKSwMBzDSHiyc5M98OXlf
8tVjQHzjN3AbmUbo8PkJlOUjIhZGOuyBVJmjAkohEwoFOWqREtc7HGCffDjwcrFp7O1MLQWvV/4S
V3IM5bNTTPDUZZ5p9PeKCZBIs1C7yoEx+7WRu16Xwfu44VX7zcyDppK59CiPAKW3WhTvvKcC1A+N
kbpX5k0yhk7R9W2Re6gG73pkRWcj0CgDPNmRrHtc43Tp4n8OFrzgMJf/e42J7KZstBJ8suMY9npX
zp5pzYEwHKNGr12ATPEVPiO9xcbbvPbGRQg3BKic764katdx0zqbGmc3i3EZjaZxeKa505pocylT
aIL+VTgi4sVPli3OcahhXrmlAyIR4r26oBaE6tojmVUBv31uM61wUQVVC5k9hR/uDN5omsZEHnj7
bK77UtSMY3o4M0dn+2DXiUEpY5eyTuQp3yOJ+zDcYsKLkSDXfSgKMxuD+BM3xgyiJbmIxeWI/nLP
3D+VGWP6DCQSQCUzamQMqCgeM8PUnSmI5FMJNeJ/wgUgBdBf8/mNuQEB3STgdtqrJ4mS9JZSuMYQ
mcmlIa+iZoK1Zle5/fjLOHSGgMEDlHiGqQcMyBcCw7VYnQpx52X0Fe2wncQHEok39YsYTaI6iP6a
q2kF1n9X1uuyayHE9Y+xuA+nrbcei8y48eUkihp8fXmbsz0IqoLBGhwBgQEtq8v2cG8YafNy7eUD
X2k08cltq3tQp3vZXg44qBoehiAkNZmYaWTX3PtIFDNs9bGUzifQ46eC8vc65GkAHZKM17LtsHUn
0rEVIY40SevxtMse+mnst7sXa+mPraG1aZewkt2fHLlS7I8GbPkG87Da7UeoPAqR4UiCrURKjeml
jRAFcD4WhQJAshxK1mtXKAOocNlYJXSWa4fTCUMALho5AKKFS66Br+9UmQ5p4ovbzwN3dQpc8gC/
XowjRn7Yab19wXVytxUlnzlpFr9Fl+0178O85IVu/tMVz6ulMdijfnf9G72HVdfnKyZ8bjBsEegv
KVdqZiq1AwMRUUoM/lG0FPWafRMGFWPle0QduL3e2K34lIUX7+8t7g6s+yuwbI4oicGqWLA5Dwe0
XcM48pCSGP0Y2Brrg0+5I22te/egFT7hsLIQRpLo06j1JlgciTZTiKHMMC2Q+ik9IU6uktds5Niu
tcVgnoi3taEHklg7o1uITSiQUB5KDIwYz2jtr4EXu2Hl6+0eYXzCF2gRxBslriIUHRV0aZrAqnO0
trm2epiMr/+Ox8pqhi6L7AiLJYYhfMgn0xi0jqY2NG7i33GFzFCHO0KvTU+9BwGfKNrW/po5qL9n
u0R9q+aqnGEVu3dGlGEcbcHoBYKnb8PgX6jK08m58FOcjjBcrMEWG/OUYdq2HfX3oSUi53Ykzlf/
wfCavm2RZsBWRGUI1gjtCY8p+mW6L+pZQOm0v8NxL+Gs1KSDyIYU9Ft9v+4XojkzG0x9utJt7fMd
mqBcDR89b5oBL5s0eTyrz8VMKi4gnt73WfE546dc2lggb9bvKvijep1WQ+Ysypt/fVohcbUotGcH
q2Kr9H3zHxyrySURbq951P1owKy9BfRvrdupBwqMW2Z6RjA2eQhsIDmTto4C1C4MNPqDHj/kWLQW
NIf/kxF/bPMZe9vkX7M3O7lJeLaFo45qFVYQu9i51OHjXpgdeNdG4cZlClHJ9M4LM5j4GCA6LlTj
sj+OO7hjQw3C9Neg21cYKBJfW/cRE44/M4v/eIM1H5Tc5DwLS4oyVTiZl44kEmBDwdk/M4nGFCGd
Gy0qffz+lZzSj660EO+/R3YWZyRh3sdRrlMHVF2gz+eeRW09H+xhutReFte/FGyibCckMdXiCHLS
wJwwIeKrZs5HUkWzYBUqMYyLutFQgRCX12ioNubZNCfvNTncQsFdbE0nTXtfHKHwgMdSgawdjYsO
S6C+BxU/tEIUJVAjmDP/dEEXHq436qWFLvUOhKTV9hWjCdZlw0ar4dEHX/wS6Kajq0sXyC24UaEn
IoNlsmuMYzJkPqcXMBJTbuPKrgPtAtqAsbKPWQhrPQq9KqaFLTtIuV21fB314T8MtXeeg1XpUDGh
2Ihvf/VknYn1GDbrgzx52Zw+VSa8CPRacv4D40hLJM6lYthU2lXcdcoEeoMIiolHegngKBmevOTn
mpHMUfbWdpwgoZTfejJoMjiAIKaze9tvPoFCdxCW3HTtQpQWWWtnLv7oo3gl9KFfKgAwkIPEO2Gj
FbE/2cf4JuD0XUb76MpYJgB3x6JABGTWLs/z0RDj1Z5/r8+qpLNtJoOJIgMGuefxlcxccLTVFJGN
3MWy3Yg3nZFde/NTru63p4/pupDUJUlZCBIpkZ5RSXIBGFZ1Atn9sWwM3pJ/Yq0McywC9MGfmPOG
rL9Z1fRnEva1aQReQO4nNWGT/RhbmmBfs72hQtQz1CP4VdzQ1RhDz1VKGVuUcP63omOD+xBbwOg+
foUCmNYzkj5cnKL4bBJikkveN4SVi6Yu3iB8sDq/FttBXD22JXNkhOZESMhyL/y8RB292bNdso7I
whUfmNYHzQStaBhriKZ39HLAg7qYJI5J5A6WCtEKkcgKsuAZw/mT6HXxWBAua/lx0a4btTro+7a7
YVh3QH2uMUB3DmVMVjtUd11/zHQLuqEEGZT80jqpKI5XNJAYAzCpLV2fUdtzZ7CItRjO719EOU8t
2A0RWZ4ctkDIm3qQaqehnANu6IwqcprWVK4O+fyO3hzbbOt0+8/q9PQpk//1OX1hsYHLVtvwJ44F
F2uhtWu3CvSkjSfSf+LHzbjPa2HczcxnPNiJ8AnikwggcOXjTKDjtpFByN0KE5ryPzNAvpJ725Oj
Bo96vdm0reX1k7588YMNi2GzBZOQSs/+kuJrwYZXEbHHXCaEIC8hSOAVv2oIDn7+MjsZNfJ4cG+W
oRnLJdQIml6/wsL7PkYYfJFkX3kVsxZOxmCX99i0zOfvBoFTg9rNEpNMJLAcREIwEeSGh/kSqms5
f+Io6nqR1HCUMQy57K+ta/ULg9Juk1mOa5pJ0hlkAIhcb5SHbPkRi1JZIGk/wpkOEqYM5DMsw06O
te74vfqmr9CH55rfbevuWGCZOp3gtFvOiCOv6bPeTnPwxe9Ttb/J85Gfl8ZtTu+Tfw6ld/UGyRf/
Ix6267bAjVFoVVykGZCi34i3ml9Zk90jN5RpVhXzfxxrkHugxce9zCRdSzG2M2PUQzTo92S+47mU
RMpXnENdNBZCfnnaxzgK63lNkcIkOuDJ6UYYNQRps6+LOPvKLMqmF7L8coOP8nr2MYjRbL6hpsv+
j9qvCpc+pRmn6qE0NWjl2u3y0w2kfvuYV0szvRU6TdFBX6iPGRKU87GptRrBXeIJv5GrEKV2A1ss
JLiv3bEdQdNDsq5YhNz7GXjMH8oK7fTyri9AX7MPGvY919LErGA7JibjM9sVddBnSw5NNs2jnXFl
vi/UbeGoqhwct2PZb1zikClwntkR620TV1uxLn16WGRf5S+u6FPPoLsFnbmmMJIW8MMHpG21cD3U
Ss9HTYX/ME+8h65e8Z5XT4vVCVo9I473nWVcThMlWNVVvKerx1xRmwqy/eBmA0NkVvsTuNzB4jjr
EJCngRgjhZ3qSLDv2rWnWHSzhWfdeOZ8dWCOMPWXCU10g3HYJFr1tOX7WjD+/awS5iSk1L9ludUx
zAoXwynS2yxoYgLrQB9aIFU08OjVf9bO5PZ/X8KxP7EmgcwqZhCMLvLAieyN7ygCF/IQsbXkDJ0I
ydmS+5i5VvYIBhOcCvu+LXPu/l/VNqYHz2vkjBy7JpKvuRMRGt2k8aDYhtRS3jV+qKQ95osehkrb
N8RF2RjowXSSlBLkhwZvux6Jv6N0VqTfWLEtq1DIlEm0wMka3LZc4f4gW0IfyhGdJwQYVROj74Ra
V0td7cgG2EeVGeZfX9uAB7Wizd/ezajVyb94uoN1komDdLro5BozOIHdXuRHJUqZq2Ti826OwwZA
WAs2SaNISCeqxg/3X+0mO8mofrPD2Lk/YAaqXihAlHzjfC3hD25hzG9pu4KnA6viv4XIAYeQNr2/
7ClMvt+rKzmxjmO3cy+tzRpUbRamGL/XXRqcgsFELdliGNzvlZXzZNGRNagcHV+N/8Vph8THV9kq
bzVA1VsR7fIx5PE6mbLVONj92rRWIag8agqwT07sZgQjIl7VeP2TZxD5FV7xSYfL7EDwK+VVvWrR
T2rpZ6nT1rDnYPYLzGAU4nLVSo1xNDHJL2456Vq5JVwF1BvxJvj2aAQdbigqGcCLuXnmGek6N4tx
fKkMJtXkCcYWnedNrBlFi7Rb4lJ96HXAShc50kxKzSyJ/0trWgtiVtMfVSLBzQIG74aQIz/hGTa+
Tj1Z4nJqKXdLhwUn2euiccqK5Z5UM5ccxJJ2F3HlWibuipwub4wy5QLeSUxQCp9b71iip/3EK4Wm
chCA3aN7tHg78OUyY5sUhJ0P+CyvxpzTwI28cDoCkBhORyjEX93wnNnNk7mY5bdU1UlxjvNR/D8d
ddsdVYcgdwRODncLbt9+lgv4ZkKKKt8DTCsCbs24gNiygd6G5hEkVZ2lHizHsbzTHwSZkLmkqkv6
QxVPpxQH6bZUjqBXqUUkbftzXmvdAp3AbWnACDHz/9oE+s3tNIhv4vG22Idg2tfYk3iqQ7ngm6v6
pL3qnbwbb4TpVlXk/X+JaDJr39srIaQG/+oRCu5yd4D5ZhD1Rb5Oq3G3UQYmYafIE8OovgTkA7G2
/xHnG/8pSK/YWyubcAqS7I/fBvP3lQO4VguBLd9YH+UzCP71PlKPcJqVbOzTkUnmMmWgWKj88ZK/
DSevvI0Zl6c7yPJgRrmz7mY9FjKHkGKHZ75VWwo+0wpYp9MxkP2ThyXGO+yUqUncfdcKdoKIA1f+
TKudSLsIUABHSQRsgTuW7JBjXF7zLg3HcZ3c8uXfc6aU4wc51opsydMp63422bemLAwxD4DJElqu
XO1JFUTiweOiXNR5isV4tnp5WluLNomDoaBVzpJq1UkTkerP+w96SHZvAkenSRNB9OthPwIlIyX5
WAMfcoLD0qXxBz3MvMzU/c4fsCags2q99ZQMCH33KTQYIR6N2uhUF5vWSfDFNHVVtbreK1ljQUGR
pJThvskt3qK/oNuJksoacVLOQkuLdEeNXVRIWj3CdUB+XxOiZ22lcVzOz2FUqsYqBt/8KbyiwRBL
ntU2qmJ8kxb4AqJh1VBMxiM4d31HvBHLzPkdijw0ayC5xY/9gZtX6QqcZqDJfsSppfqsG+FKP8OV
E4ezh6RPkCCFliuOwW1jjVyahThvdvoLuhXvwKQ3gQpTbZ2Zq95OQWl2zwrQ1NLwul6NA4vJqGnM
WW6lh4Qu1CDSWMWaLYBwQMabWq+9j5RORmpY9lB2Jpn6n9Znlm4nr506TvfiEHA7yseYrOMc9B6U
YCf6cZg6PMNz4KObNCCO2o92c5NT60MDJf/v0maWFcrsViC63IhacGsbeXdX+fXYeaH0gepe88go
Jt5vWEA+7WQAaoD9sieAT/r+Kg85TdnQLHGeLWAAgbvC+bZaOt74IrfpEr4MsTIoIn41HlbP38vs
NsOZem0I6N3HD8OLKeIP50NxYzo7UaH4lqmyr3KeaA/noTl1lDAOb0/Ko2eXi65w3Efmdro3pBDX
RR0qvuKT3sTfCatk6Aq2v9lTxuUJQpbBDIDgCr6U9b4Og+VACyOJ73HVtFVZJ0iFKLDGQYr/pZMx
n/gaTKSUEd2KMrzn/vl+U4Wk4rAIDDTzJmlyZqqmFUSDjIXcEeY7iKA8iqBS2K8kDNdddHCrR0rL
OY5F8MxGbPsL8/wxfAjQJ5PjqzmyflQYOTsVwBXEFowUHCqe0KWm6OI+YbC/1BEh7nuKYWzFtEq5
UhMVu2qe9Nx/BYgQ/8Fz43nekSUfZ8u2vOVl4HgpS3yjrJSsFFlxp8OBcmhBE2fZzUUTd8Fkk+fW
WDKE6l4p2J7CRVP8YwK8aCCFVTx1bbkWR4x+hwNObxlXWnRF3t8ZAJPWn/D564mn3XNWlh9UoVxL
vsVCDGhNWxyfOIGZEYP7pHrL+LuOtzwIPGhCVSiGYZ0f4nz2XcJG7JrHQ2DU7tv1EMwB5AnbPHJD
6ea/Nfu6Wazifgz1PYA0CXS7+rCpGTmd4bmS9pLbEaVS4UZ3ZvVKjPaakXXPJB6f1DjloSebT0Iz
mBqKNhA0wQ1MdWDm3WN5X+hq7tq+DlBthk6CR5gUM69RR327Qlw40nqzRTybkpSaONbhMD2oLhOz
bnYHZvEiqz7EG2qpJytTwsAgjEWvCBxP0d5PwCCKL9ECHEpRpAJyFSdyU86euVdNV+fMcAgRTf/v
xGJVt682Jpi5ImfGhU/TB42hbz9T7G6W7AkKoOswJbUHhFwZnSZa0pAr852bZ3zuiqhDKLAQJibZ
5U9oFZy1yNcNQkldEu0GVUWzy2cPMd1RGUAK+ty1J17QSZ9u0ZSrG1v7pf5bKTK8SnpyoKk9Vg/a
Pg39sJiBV1XfiIaltcKTF7bPeoDeps0yAEvs74mTnIa/7f6+SJpasvSCym9lOrehfZupnkOYIAh6
RJbxMWY0yjytI1zXgTRpRd8CjN5i+Rm5RisQRrUFqCxSDu+tvhWe2cV6V2UrRdtnHEUkt1+vyg9w
cTzZyf0HULsU4ogQxsNt2YULJcO1XtHWypD3nw6/7MxiH0Kh9PvmQNb6NyVC+DekZ0ccwV8abb6I
QaSigREqS9fo6Pr5cf3/TSlIkjtTHdzqDL7JbS03EnQbPleDqmrww6GqdoxyCYmFyag7PCDk7EfQ
Cn6MS5L0N0qRos2T9bWBooH4grxyBcwNszS8FtO4VZwymlLOshOrY0H6iTQ2HJlmzMAtmyU/2IdJ
u6zj4XbREuQokNR3DpLcAqTpZ9YUiBYsworAwI7MC0upTLIIvtJ41zRMUL1+cDEOztii3jSioon8
nIbWqc5efoIpVioDWEoInqEOgjXWc/CGoHAGKJxqepyuE/BaJS8NQTIdYhjBFR+RyJv0h0uxPfuC
polsyqtf8AWfG0ckPHfE/AmcRLciQdcBLdDe1SVZbE+ABytoRFfcU9Dqlhu901OJ/VgDoSI9x+gM
yJJMZBYZ9eLx+tiHVR4XhFluCBSBW6FZzRVpX9pXXdixR/rMOYQhz+EjdaiEiosR+ne4bJaDuKws
JEVGyEKd1ePe/m4H8+JNGUVAwMN3uk/dWjnfk4bIakPephjSrY0oiwsKaOIK0UMywJWgSChQcqCj
10NoX9+nPqUZ1/MH1euBYYptexALoj/NdTaGcmm0R2yYOQqpH/QBMph8Y3mavA8AwWgrxDVDEVRW
xnvv+Qig0QHftA892/9Emubo7yzuvPT3dMTZ/vnDlDW+sRUD4K5Ju8jBG7M6liAKlRBgndVUO0Sj
EBc+3JgSCD1lpUIBt3CPVPB+vywHbDnA+Tax7Vxgmv7DT+400FnRfEYrXUJ2YeCOT9ogJGpXWOZJ
NRWjAaE8I68jbVAG1YXk5G/kax2XldXF6RDjyll6NdcFjNVHR27vVV99ZkDHcWYgJyHCEFDvCgQL
8jnJcpm8XfDIJuL0mPmbSxXsy5Wt5ky38mL6rwg+tTMsLfgRjrf7jHwCMQIsVuG+SYYi7ZQztgJo
HmVsM4X5Igl+5wofDa/HARa5FtR9o7Zhc86Txr3zRjIcuc+1f9cgjo9Kv6UWZuDVieh60YfXa8UD
Ko+juqVHqY5xVia5wOfwti5lsQQLlQv9TjIQNp1uoP8KLHrQ3PfF5wC5C6eMOOi0x4dfHeKiZANu
atg+n467tnpZ75/SukwIEVtA7qgFDESxrST8ofUTI/yD+ecxRA8FJQ2wYdy8xEdReW5YgLd+2EEG
/WKs1Yq19gAHfWbijo6mNvt8kPyUH3yGz6ZK978/JoI8kMzoL0hWlGuLXDM7zSf9Qzhs6WYy4hEl
7U/VSnVgjRyTDNM/85rXzQBITgLIp5iGam6RNtzUYEDsgfesS4MdjiZa16ZxdWdT9Eeely/TI1/P
f09Ui2H9DC4sm4IkaZBhNzB1b+/+nPwVEKj6i3rWa/063ySpPeA4FHeR9PcKGks50KYEv++QshzA
dLe+JmSTQDw7U7hZX7w+o3QVcVQfSMBAmWjmzUiwvFQEncQqfG3+rBYZuNi/MSS7yhwRXcc1SPn6
5hpUgsU9EgnVLXjG7FvsTq3LE1A6KsqHR6+csmEt5UvrPluTkh5A49pEZlZoCXreib/4ECtRVr9E
IuvU8nwyacGzihMenyXvBTTVdhEpYZoeOBd5LnI/kgaxHIkQZnQDL/tZfSFlfMR4iyulCjif15Aq
B6h2icrhRZ2KcIlEOvHtCxSktiGOdMisC6DOT720Q6hgSTggjqdILPqeHbhu/hA5LPHw3HQWAxfZ
jPdKpTfmT3GGd/u0QpFl01UGer2anIcWI68skZJyYU/6Um5AtjxXVl8vEPNmlzG6ImkriIvY4cws
RXPn+1+Iw8dsUluRxva4xT6o5BgpJqQp9CBzYMdNu8qE66FWgI2tU5WR5lWrXH1FUoE2scjwUwwf
7kXPGckGODhBUB0xrFhglXSmFi4d+tFQZrGFWFkMYS/0LcLZ5DY10GhSh3F46Lq1JaN4OcnNp+vq
LNQTVRbrLa9wPTJE/xMAhWgJYyC+BKKTIskaccR3ymRzAGturdKGY+1RsvOB8pzSH96lELEryMHz
p0htaMMwQWOsiiQiy4/x0isI9bLar3/L/G3I4+xwYd9TyH1ezYPOwegwy2B+8gCN28mbUYKo86n9
qeOWG1l3BgAVMAchy7Y2J8ZQFM25ZGEByIHQkiUgaelQ9HM48BLr+IiyXGMehzpg1v887O/H9wVS
Ng9HTX7zmFlALgAj06wWl5jqSClALNzfVs1UeQY7qgWw3g+/UfUbL9odQLuZqijrM0Mg+Qs5//XS
wQAusHVJzdSy59MY92oiNj4rqrrgzECQlf5EqyPATjI5x95m14Lg/r1PnlJQDfT/8z7dIiTQEyNB
0YXxb9R0LBtnUjs9EXtPj1l7w0EiW7xpny/W2QJvUHFjgogw5ix9NiduqTFgt1cpEAST8hE9y9+c
PbDr+S58/86tW9j35Pu6qYmtuV6VkCfkpxSGrS100dLZIuop9m86lyZHrKpWcwdhLQ95y5mm1E0g
cSd9ih3clnrpCzf3n5OsQKApPGJQUmboLTlsrdutvvZN2GmRGIRbmFeoljzv2HC0c3IdUMbaXZE+
pujG+H3CfDdUq3sZI/GChokfh9FMMl3yiT/MV/2ArGnSKfs/icWPVd6WZp3pXmkMoVF+tEk7ZgLc
J6cB3uzzJDHGjJ0pymwlPszrV0uZE0/jh8QjNGLNMqkWWXxpXyABeKVcLBTnbQGahNDoF4CeI3oJ
OBjSCiU6L/5PSd2wz9fSRV/pgrEc7/waTcrP/nuh+BWdId+6IKY0HXV0SrvpzJBR4pfkGg4HabYd
C2PYfbZ3rAj6WjEtugti5KpjZ1/wGpUWtZPGNHmkEqcelGqyWJN7fos8snhBjFCOvcacIi7NWiO/
/rr7JGsbN7K6kpU6xbhpw9Azd8gkvYhFxrW0JKo1f/qWj4UOzkj6cYAyMMDQFW2h8rEDsawWM5hj
W9uhl9nFX5Vc2a93ZkATTRcbte6Z26zTSJ+JmlWLSQzEaCwFkIdKggPPWMQUT6tdRf0cgUBokTse
s4vbAmXDsg34eAWNZCb+dzW5fy0CEjl5B5P9Ajv09ZH+FvFCgT3SlDfSbaSxQppdMOLsu6qblZFM
uhfpo5yNwYozQvCka1rLIJikq8PeqEf76YjkSH5MmlIP2SFASw96+oBnaeR52HzxSZwBX+kOxQvO
yO3gO+z6fewSvwle02lTdosC7Q1pwX3zbrJyhGs6bsfwr4RM9LSl3ELCiKZB0fbp0aJ4HQZSk4ae
bTEwrn36qY9CdvZT5XkXWKHBKiLBpAma1wL48e1jnoeGGu5k7Bo1jlnaFv8R6NVXzG2laxNamwX+
2BZuswC6NloftB232TLL+CcboqNiNm48VFAK4d6mo89Zlujfme7N4GjbmCkP17zbp8mmTZ5YB0tA
glc8N0sdoNzJ21WKBUEF4jfTrwC6O638g8h7pbjPMv8KoJdUUpsXisc5jUj+YylM2nuSQn8geahJ
NuZTA8bdDZrjBvy2KPInQ79GT7xf/9zrJE+oBb/6eXxM+ELYYaqRXR9RNmqsJHOya4c3rDAX7p0D
5SvBBplJgtthUjfiGJB+Hu+sJ/ruVmD4OvHbCO7hI6rPE6rEeERLWL63NWgnNQA8sOyehtAZKHKX
1UtECnw3gDYs3HMwcSLfyxtQ4MnbQD1A6KWVT51FrVztUanVO8fzHsig1IBvIPUBGwhJ08bPzeIu
74tj4n3Fuam/8OjR7iLTilZ3oA7ZzNikiy9Yq2k4AfDF2t9rhHaYvZLcI4HEPDTQ2CcJJqBv4cs2
IWxyz/31U/MCI00U6VP76IxdlPnUBA9EOLBz2XsZ9rJYOUfrrvzn3DbjSrykaxlluEBbRCaOnWfA
535Abg9jNLNn4PqTKRni57S6Ye/Dba4GbxeqhA6qYHx3fkou7iw34UnNSbsN0OPczNhEE+DwqgHM
UwIzvD9fhSY7Oy6tI0utyxjYGzDGWzRkmaLMddtONmFdN3ZNLe3UokKTBMXA6A8Rwciv2uhikxIr
sGzs64XDbkkP9zA0g4ydyNvT6HoZL/KE1zW0FsY9BJoEdZHtg/5LyVkNiVdtZgNlFdKS88weN+ql
XC7NMYFJ+8Jjh7gJOadeSwk68IKRF6JnfMoAXmdI68xzdhMo0ogt6trVQHUNb9JbUFCkGhbnJQUX
TPPenLcnWiIyDJ/dvFiGPdRTmEGVH44Xqvm41ciqRQM2UPPlPRq9G/D2HULk7HtwG35p68yOzbEQ
/gFQBaA7qK6f3shtSQqbZ6UifVzt3Ekf2V2ZjrZ2LuhKd8llDUxG1rQRlN02yMxxlxNuwn+zBRaw
c7zpXuke1DTwgotlDlw+aPbf1dLmliOVtWwzYmvIZQgqQm9ogs5+tR/7SNps1kgadIDWnjH8aZt0
Vc84EQYrR3tZvFviIn/D0QmIfD7+nXwea9Nv6zG61Uv/SSGhDWkhLRDxwQix7XOhmEr749pWWIQ4
JI3T0T68nSGi5Dvi9D71lfULcbNUMqEmlUdRjAmgtMigh0uMYeKOceOwtSPRk1rrrrVmvEtZWaqu
4T47iSNyx1xWeYdWYZ39PY3CDnxL/gWT2GAeUn4CIlpXxNBSvSBTKynREAUQjguVCdS1LA8O1PHs
v0lWoYz/j53uzzQ8ikYnVUMj3+Eee2d2eK7YOVOU5YwH8Dni0d5CsQaF0sxVrzQEXs3XYvxRn5ZW
t+1urJmnPCfnzOWLGAN2UBh97kCXXVEmLi9OkgMOxUJQujbitSi9VitG81wfZFUThOxsuFC7sbYI
h5jTPNi6i6nuTUakNii3xjSveT9xaLC3RdJA6b+mtuws2nKy7too4pfzQuzlavSpbjppjHa+/Dns
vXOEOrVjmIzIINchre9tqnFsO9261Bff/Bj5fhLUXtzzbY2QbVymqB1PnbZtvT/bxn4G9c/WR+E2
/ga7KZzeuVrmD+2Hp+5W15VsZGusaGpY2NfVWTrE3D+8LuJc4BcgjftCD/3pHFh2/tc6RYgAxSnw
bbGhFfHNV+koUQ95bf+PkZ2LaWD1/hgLBv25K6oifa+Tx3P034ME2Wh/rTO12C2xP5/sZ4gpvU7h
OfZcuJ7+ZbxQJJBQ+86A1Qzm83183FZHnONpU8bjXtGDXN+fMqOeMYkw+sQ+Zz9UOXdKBqO/mn54
lz9ICJgjrQgrnOFzwqxaZjpY6anp/vL56p6lZECUr5sndRSDg3WRN3qYr9IjfDi5FR0EWyXTk5/W
QEJMSw40fWR09XNleG5Hi7bHJwcRHflmj/kENCxRb085LlfAw+B2gYi5qPZZU34VjQ0B1sTqvpc+
679TkUfcOwCZe3O4a7Lqn0P9YgeBkdtQL7Tyd+cLtCVGXjJwoljJBFOImPgD3/CxtvpdmKQdlHI4
sko/xbyVCSCMkMhkPy/WW7ypSMnFf8qTfcmGRHaiBmb9++EIfAIiJD+el8gwIj/AWSsIsrirZfyf
pzllw95soATwB2tjgFSibr/D2jrAbPUvvYQXt7THPySpRMuHO3q0eVYXjKwwv51Y+mbTwMwssBex
f5bCRfObZyLs7PbwMzcr5JVuXji71lsZIa8g4tG/7/HvCetMc62dgxbhAyYjMc1Iuy2GLheI9pUb
Z7UH8ga/8L4dONQ+gPVbn0XkCe0hobF8inlstEndEUoEbSdsc8rcSqEsArTNE3cuUwtbPOBhYRfY
0qdqt0vzXLTboc2RMrkPALpdOuKDaw/kZeZEcV7Njj5pXlG14exndfa/jPT0HstbmynESrKGFJzk
Fs0351M1HyZY3+5hXVSoo98ps6VV6rOMgww7MxgJyWUEpWFn6MHjx7gdC7zfDjvqrulJpIDBF5HC
79vQ0A80kiYleacVBYRYpeZ1Qq/zWIQeJQHIB2eiNU+jtkhpFqe3Jgp6UKeH2mzmVs+es1pIZ41q
NXIMcXEwWvfjvZr1/zUerS5RC4Y2tCeoH35qM2q1dVyExPcDvX58HiPRLKIs75Kk++eXnIyqhk+0
/2fh4Xu29sqnLLQ7JyuSQsOMcc019ZHOjcvmXVL9rTKR6pBLzMHPhzBqdkVZMKKXqFVPziRHGDHD
p/8vHCtD2d3FXWKNYySZfJgFW/G3O7g5f+YNIjX/UdlpsAZKkDC1rhnexiqPRpikDZlDsCvVG739
sc+XwcBb9OT5DbV7ceIPPtG0HCypEH5X50dOv12FgVkF3kS3vhzy7kE4c1xPQKIdw/zcZWnhzxQq
oTshwxQ1slR3EPM5ItLTAsAReRT1Zg+WhF5hHoO8kY5/9vcVal8sbYZRcEjlWSrj9N3BIjJo7syb
re6hMay+f3FyAaj1wz8zPGsAbIqtMoM+DEwHSCXONa1uQ2fFS5U0fyX9l8tf6Po7GNAKNhFhId8X
SFPQp9CP0qrNPFmcwq5m3HO/8fDD3NtyU5fzUneMG1KuGujEhizfRVulWLxil+CMXygDnfc0EPBF
/+Z/+zllLXsuAyH7jvhCId5zFunATPWLlDr41BxDH5uQF4OaU/u0xl0DepcfLxn///4WO6EpDL//
dslEX4NpkNgl0On1ux5LRt6tUJlkgGhaqmhm4GDKvpthdLKdzldUUgJzLBKgnD9Kyxg3mo6V1nHt
mqQ+ePlxOTgtdi8yrn6+tTNDEtmW8E+PCZB0TPP/IcYgbhiXbt5soaErRonMo+wqkE98mhWSlvrd
fUC89Epn0qwjDQ1a16NVsuJK3G6lst+218Cg1NIv+NCHTE+qpx/0jaMg6vITeMOECsoBvKt2yK6c
1M+OnShUDKZRUOiiwhw6aQmdUVm1RXLId3aQirOOxWk/yXVq0Wy+Ot9xpmwWWmjg8gYOnKM3D0aG
wJJ3KEi0fn/alkqPIAR1HDUZglD96ZREvnwzjX9pcWo+z03atJlKV9Keyx1n4vPrlV+kiTVCsoGl
BCFymRkIW6Gx0JICdCGcLlHTwqesUPgkZGrPbthanJhlFEPCwa5Rhy6isvJfkjAlpL3DdCXcAqz8
SXV6RvZ8jqAEV6d/SsEhf7/Hd2wbwa/+XJ+aH74wd7JrpkA5xexVnnwAOhNJf/4aGEPBp705oFsS
xYn+8K68rWLkCyWOjH4jKY4AulsOwo50GVT8EQii/tw/whIMGHMoCKXDdW9A8CAtg7y7k3i0nDoe
2KHGt8CdZTFST3G3mZK0BRImhr5z+Qc5RQ+zV9b6zfIlr21/fCIkaxokYMjffAEAkMgLs0bfpZY1
8CSt7NjsiW4qb8/2uLuy6TBuxy5NQrRP+O9QTodwrpaLjMnDLAzdWNOCpr9aofkWB6L++wzgp2d8
RS4kTUtAFnmJ1cSTdB9KoBPMF5xG0ut9/WG91Z4j/i/W2Bxbau9Vos8oTcx4BXKO9dtdSt49M5m2
mrmr08oFoZvWWhCzqImi26lw6ZEK4BKPFGMVB6HsXCY/h1ahY/NsJr5AqNTdG0FmwUCK59iPQfPi
dXVzakUlcZBlDDNQH33wkteglxJZ1Foytq4s4lw7RrLKr+sApCIDX4a8OehCGF7gzSgKaw1sdc9B
BWQIDhiIAhVQA8gO+jQSBVAF+Yup1LphSz5BJiCBofnZNUMnrOEv7YBPZE/lckAU07y1VjMOJogs
ZT3HjJuNtjVavVaapP9/zH4rjYA2hDaTuQvULTFBoylbR91QgDK4US5lFRMGCrWb4TcLOe5arjf4
cYj2Jm7EsdDIVYEueH5Wq72l4mPnk/VdkO5hVr3z48HZZM2bVNwvk8kbYEQhi8u6tdldqmsEc8JQ
JAT+3q0YpYtm7uUgUxmG2ug9BOt5XpD7z4XiNm9NCqyrMg39edQbBRvo09OkADOiErxj1j3uL2ml
MRmdxxC4TYdAG2rPpcyzAqsRDzVHTdaU6Ced2XKHwHuW1NG0MSfIWT2OFx5ye1PXlLOE0puMFuSa
DFEqkbi05VC1KiYJhbmFTRNcNnCryyvDBL2bTCR66c9/WeBzrjO6W9ptoj7dI+D6snuGmXoeyWFn
IN0sSJGHqzSUWIimv/jRZ1kdcEePMrpMSv046GqUv0ztIYhuQxudPK9PSX5sQffc9phrdYvhUlUh
9mZuxhyPm0G/L1P/UQSb2ZsedxezLuhleuiAf5tJn5Q5ELDL62UZZZlGYLae9XULxdM3YZ8xSrNc
z0Pz+RzRe/eYhQZfxp2D7b0gvIS+Kp78FMfP7Z6TAThlPOk5gN2YdJSDIUQNWyh83IS8tsM6/kRM
7RGqoIL/fmj3g6VINSs9fjXtER3a0flGoyYkmZHOT82W8rl5QspgWcfIz/NBrAf/UAP7jUvHhAVO
qz+tmORLoTbhmOiq6rD9lipqZ0G1E+xnYv/kR8Ok+7TW0gJl6PHxT+m1IYS+3KYkZK0vOJLfNmu/
mfnrVkLU5sZ2QSNsaVX3+8ivXSnTTV4m9qFAxo8nh+qMWx9VViEvKd6THb9HIpHIWrDNN7Fn1Awf
a4SWPvZqNb4v7pLSzoBQCZ0XBnaRDJe81hq/JKy91ZUo5DIccUn/pj8GWkFnkThcaaW6jdiJB5VR
FVZRBCYfFZ0OXrkHjew3CRPM/oRaV7AAXiOPfF3nXBJAGuZJ8jIS48qo/EOsZEA5BF5aC653JTTY
nI+afQlLf/rjohGPQORs9DgMQeCFkLDzuYbt3rpdkTFic9a0G3/w+T70IYMDOAOP2ZyKn45EcuUt
wlWh63FWytCCZvBhR+7KEZgp0BAs9pVFrp7LltO+j4Bz/lytG4PnCqI1acPRWGxKwxGqg5ILzEU2
8HFXHRAZBRvEy/y/Sfuk87FkAsin4DKqVWJkHeLVEqOFwcGvzLJWZ/RxeBtbGAfVJMP+Bh5k/4YZ
HaDgVBewX/xb326V40I/5Hqq/8ZSllTDxLVileLUHPPHZIdFLYCJrG15PO7V9/xqYFNvP9yBQhJT
3pTxR1Psyki5pH5jN7CJxxl/UVs+alBFMJMWTOeqojs/4kHmi0dKXzrKNJ0DeGRfN6NlTtj3AScw
bqFNCAfuqX1acdofsEFzyF3S7S3iqyCRPpdGSXvTRvXfbqJf1U5ewlbuqBlkkeutMijBPIIbXvPg
mu+RkWqiaZQ/jI1DtSva8cRdi6Lmho7AWJ2cAT+muAo0GUau7SLKtEJzzSghFHhHrKzQvgDv6t9V
DFHklRYeCIWjANRV2AJdfBUgc/ky5Z7Fap1MYDOP+msm+lZI9N7V8NG1CZt76q6nLSBK6r+9pmr6
9bCBB34jfxnQODqjA4ORmzdRSFCs4siFviMz5IbTeV/+CrYCcl8FfnLu50WyYWUVJScBKyMJ0wrh
K57gBFkHr/BRsHqGO4oR2411hJ8pAbMiPIAf11yT0232AomTVPiJTk7zkThmrWACWPl0XAQLwGWh
Dei/oqQ5m72+lynf0Yw9xlqOonYYug9RSYvVNfMrJYAEdfz0OkP/0bdkBMOl7O1CS9Zr4l2KYKPh
I3+bXHrvnWXTG9czSIjurqgAO64xTPvgAPDe5VdUWrPWNO+NWLMtlnktvPhGuf7rb61NHp1RhGyd
iEWnq/3o6Qog2Ndo5oH/bjqjQB8RWlsvP7hxaZHCtWZminnt+/eQgTkCTHdVReAw/qiugIq0loTK
4pu6zjlDtvGrp3T2WKK+SR6UEZE7MdYr7ind671u6nhFn9n5EDWm0sJsDSvqkEUVo/ZI9/LHgIVD
VHBB/pmIrJbetYMLRQ6yaKKh8J94N7lRrW65fJCklqIt/6Mer9a1f/OVeCnImv9N9zU1rn5GG0kM
kPEbBhkjxWhHBmFS3pskeNJqCcuF+fgaA6dZQi5kgtCGryj6RGYxWLVErk2mIhdErvbDPOr/ShFb
UPT/y6Pavv9UilAbtJ8uJpGJtcYX8aXjYx3bpkqKmeO/4lFUiqj5aFrU1cKlFlGVetqz+6oxVM6w
HDEF/6KCVYNP5SXfpED3c6yZyGoBSd2Gm5UYg1JrwOUxgmuE8DN0DqoRRxK/n1RKLq9eiP7BIaNo
PKbDKpr3xqb8YhJV5xMtsI2uSZF48kSqsuzeTqGD0JwIL7QlnQvXH8I19HuK7NohAzwzlxSbvwH1
BQJPdQj8d4+lcf3lCeOB2vbq06hlpm9pSjMwSvP8D0iGqfGGmrLMtINJNGVHvnzrkdnL+RyrsleP
0e/BaimVHLcjJqacEA78W1i6EMP8lYHXKrNF5NEqK/mVfN9vMFWg1aFaLVMYl/Peh6qECMBwkp7v
A4HI/UHQHej1goAhUVN3oh8URsHFDG7lyVxjCSiVWHp+ZgJam5K6mq3dLU709BeB7izwrEXh2WNq
A5hIvq030vjem+DxWc4h4SsyOrb204vrStDDiyWlxMX6KfNrc/+W0nku7BGbZA/BTtjSe5/6X+92
4goQ6GZj+nx8lw5mHqdlJNYXXQGHGqA72oqqlLRhpXkjoCPURrutRvHGWf2ApHtBJC2SmqhMDEXz
Y9pjYfmjo+9rBefzBUhbRpfkk7fGnpAarVjFxroLfbciJ6uZ0Yipnswv6aPCRq82flMxO/1Ynen3
90nmfaIgy4lD53tOrzOFS97bA61vfUyHgzoz2/USKU4Q1kSuZCK80MzVZ1uqrXchCzE7LrSwzP4r
3oAaWZTEUlghuTDEVPOHIlb8gdStjHZx6RGQ+Zqkyq0qiuMUfGxpE460HZrBTHnOy3ERsus/C1gx
x2KjT+M5TevczdJ98svbLsJ4DFsn8jQlcM9npZ1s3RhE1xwTJae37SchoDHqLBK40pBLWC7S5oGJ
z+PgjfwQAwpW2ilY5kj20dLYE+fXJkFfadcJh20ppAMDu7wuWaop4IXo/n9hOuFw71IcbHiqWnce
POXPh+Rio3MqJgSz+bGzgcqF00Ab0FFi1MvVZnC3AQmD9ZtgRpeSMf1B5DAqUPjLVsQ9Y7psXhYA
aru237vxnqmlqdlDzhao/M7Vgih7z9nK83W8eV8q5HSWZsjpi8k3UXN9kVsRHsRHakt9mO8njIxa
WE8/sadvhKUZEfPiTSpVVnuZhMPhXPuf/7IQzbW5XIp6vMb5feJuNFqn4Fncv9iJTRMUMO1lt491
224rZC43yU7e5LSR7at5R67Kx4v/2aGlPPYEZXWQJ/7PCyFeW2Na4Av+eY1MSK7bpKqzSzb4D8qL
sB+YDs7UojYZc4XexKkfGtI2wVQOay8PoqtkxBeGeyNsU/prsX0PofMyZcVgDm/14s4rkk3t+lLI
WFFK2NRVJDu7A0jGnEKqX6qDg8YcJcn2+TmfsOa7vaTLQKgg0yx5V1/LRYFNsyLfGc2BGcMIfJNY
lThpVIOogPUzZlB5mQQRRf2HB0bxctENGXMKszcMaFKZIstiXshz4cIAf+wKJ0lQClHgBTqFlhPi
5uyv1iW6JCNGHFAdpgpZ/dwE6fhTWG6xt1pATIEHGGFoUbi46kmkfqFD61AY1X8a+YIh7w48Cidl
WbQrKz6AUeugrm/5SbA43x4++kJ1Qqx3G8HXTxn8Zmf60XeW8/XzSs3K16xn84JovskX+kMy2Lhv
mgD14N/D1Yis10fErQmtHhajpl0c4uqmbTArGvk/lD7tvOwvDCd7M0R1eeQJEBDXVIVWnj3kZt9H
nqLJYqYVKFYFt3RUqcpwIn0rxJnFYnEBUmLMEq3ztrjvFaxIzZKW9oNgiGC7J933mdUYXHBRlfMA
H93Y398pH344ai/TxjJeEX3vz7dMVAB+kAbrhP0QS5f8xSCj4vAf9uYt52wggJmqpbkQID3fe62u
EgBg2yTywz1SgaN2gD7mRam27vzn9O571ncHXvl5BG6GIHgZCLazhgKRHnHjNEQ8dIgheJSxBxh8
j4iVJYY4E6Kdy/UJWpirZdoAHDzO51mCp38zVW/WcEyUtt34Zwe2rHLVDASMtglUvH9koWeH9tWl
Kaoi+CNI1RDm04K6yTWnFEj8odOgPJhhUeLTsYONyQAMdcIzUaSuibpdnl8twx5TisXJVp12LQ8z
3+y4kaZG5dbuZmiRjIL1CtTioAr/Evyu8LmjT+8Vu4/lU4PTVuMWq9+islxzDAyY2wZlgXacYceW
azTGECdplQEHniMpYDk3zHvd8/1P7zP8+rFyiU8kC2hrCnsQhhXH9bJCCA/xv2uS3tEhoh4fbdFG
UgfLp5+TM1UMcDUTDTtLK/46uPivBucpawblwq22K9QZqIU7gbl1WgdZ7qaXLsJP0s99skiF/pD4
oCU8F9sxRk5nIYd7T6wiHZiDXdDHI7teNkS4X/GEPgpiC7/yopoZ4nxexZzRpb5Xl4YC26YDQTw7
e5GJaIQKt/57O0BLjupyjov9noXNPtr/sS6YpktNCghecID0mEGHjHK83u9PNAKwyaGmVBpD4HcV
3NT8ZKbGaJaMwlY+H8riZ0xy6C0eaINP3gdjM/vysK3jmXvaIn+ldxRenhTU0eCTwEmWR+n3PnlV
DIvkXOatrKT2FnryJn1Tp/hZlnBPce4blkPSyXGR0mhNI4u8MANK/VRc7u414ugf9/ZmMy9xW4uU
5/WGyh1D0FifpynvTeWw7vKN91jshEog+3Ep86XuV/1O0PvhYYGamE9BZpTlTvQuc85bbqPTiKTB
JStoWSg117oPM62rvPDENqrVcKGcTaWyg6uhaeIXkPKY4WL7BgPdvNw4+Ed8G+TLf7oXdekBSGQ/
7Gk1ZI6RBSUQO/eflXGr3dpn7/fHBnwbjfl1DCQWHvoMk30ouICM5tmP65AXyHQs4J2XocvjDtgq
hJN4JSEGu8bbbGUZp3JZvtOcMxmRycZWN0q5dBviM2EzNknPUnQvAkZAkjfLupMKAHZ8iNSFbCfC
+3Xn5lT9F3FSGSJafkGkCV6zSBktbCSF0/KwZZwfSzEdWgHa0BUnvHWqdpERK2gzy708G5IKinLk
4rW76WTL+Ac8yPZ6ulokYSSH4UrUCkpF4eDNb3k2ARSS68uvzFAPElrEqsecQgtCOShDhwvgUfuQ
BBDOv4K2CWX524zMfb19WOFDyk2HGN9yiY44yDNdyYna3zSxTrswwbA4v3iVC0hnepXBtJsINZ22
A77oGR1T+dJF8s3j7+Z3NZBytxc2Xus5q3MNOvmthR6Xp6YotmWVs+5CEpEkSHXiNklB9O3FTtHD
AKScA4Xf6y2kPr5yQ+XQ7f4gf4uA4BqfZQFyohhZ40TUSmnqM0idZIGa/o+s5QWYjnzSXEVrM3fh
0+7QOsOYr/Yb4NF4dBfhxV35jRjca8i7owq3kiUrP+zfblEgmp+BJiAuc8MCynxc1WKLhOg8MvbU
gkOXfiwEPwucetkgbMGbi6/pCcvInK5e3DaSmDHwHmPNxwyVQFvkFAnMgn/isGU4/EhpdE7CPbP2
TdwsqijUhL6H2Bt3wHNr0P5yTknV4VW0WDsxt4B9j9c+1vUcKQrjUeRgUpzr0wJqq4u0SEa1za68
XAOrtmgh/+pRB5aNepDQQ5Z7Vd2w6HgWA1JMUI8df7+MM16uLpPJWPhGQUHJEfhOtcVXOddsOKWK
5mCxfesbLwaI0YrF4sW3PFox2aVqJbTsZ8Y7nFWsm2IIJWdXyhUKayt6AY1Gg8XqI0Nmggqfp6HI
sFNjsCX9O9LTeDlh8C20iiWw7utrJN6d04RUnI+fiQOcULanPzinXE7Rxai0IO9O6uUPxEKzyWFv
aTK2smNXldarQeu4237QBLeabBX1fxfwgFInUu/EYLH5aMP6P6AkhEbWmbbe2MPMkZzxdP8QoWF7
jgDpftoy/K8cONhiNbatcoud1zKJhyvVpnmY3pAl7rf108Frij3ufwZNf1jFKzip9v8xhVvjI4qg
18oLFD7zTIj8yFxzfNwn/YpDQkmTclLrj8Cl4g9QpzLUH2Nqa/Go+L+rwTtbdxC+JHXyOpHVfR8A
RnmESwh546DFGKJDZkUghc1JNH9v19zpYdm4kHpAN0RyMXyIK0bhPC0wryseYBsLuKMg6a1zEdU0
MM+0TesSHo/PWzSRXfH9psHBnaY1/zHzfYSvHvNm62wHO/Hv5oTqWi2eYGa+HsXRYYAVWI9aSvDg
vfhr47LrdCslyPKl17xPQO16c3eCLaTdVwk4OTADb1YHOXopfSVns/hkt82pVaS9jhjkeAlR4BQl
Tt8TDHsXlN+ncgjp7KYhqwZL5BDF9xB4o9MlcWqUM+3Wuh3lMgY9u6Ou7+XcCAysSWByRP/HKVHd
MkRRUNBsWlohIE66Od7L8TjL3zLMsl4+5bat/ay+4zW+/TvS16XL4oA9NbfILDEXfByHPSYT5JXi
cDekjVC3klg0EgDZvV21t77mhAVBrP9/D4sBSIVEfZ/EdEzvevKwXv5f1jBCOqPXAw4gBIe9U7XF
w5n6X0ksLNkfhGy7MxqSqOHww86fiJxAHMKhKCo/YVc57Lx7WiRhYPl1gOpCfrRGJUPvRaIF3TlF
BBLUHlNpj5BLleE8xnqGDvPC2sdaiJi4/FAn3cxzzWTPpc6aaImq4urKjIkNbA3urN5vS6TyU7Pl
hDxfmyMS7f/kxbIFufLSVGgqmXjSZ2ut495/NO+TGVCyx9fy5SRdgJrNTPqfABPZrHuLB+Yg/eno
YI3KWBi4GljVTpf6AbCAbKwGfHUa6v4UofNrqOCBKH58rLxwqDZDmebsZVA1y8Ao/0vqUCUligpl
wRoZHNBzBfjfRLayhYdmQrQB1PV1S/CRMMgn25QXnrt+JCewMLYQYAN5ZHO5fRSd8B3o08exlHzg
xW62fU0+hYOkl9dIqoP1BYhdXxr9Wh4TOiLbLKnACXUQj24ZkcVokxLPPMTKc4kcf+Q0XeAtKlh0
Ejz8iLaLNCFH5071uwdYHBEAAuegqpN7vgfLgAH6yefh6g+rmr4twZqsgWGOrSYmURwaJw6U6swT
Dg/z2mP/dfRIinQWK5pp1k0ZsqkdVnu3rZrqak87IjNsEVfCrhpgo8YjRYyeQgIIl8tjypEDnoUa
kWp+8rGabbfhfzGKYgs2OmO2+G7hz1K64pM4xcH0HDdBlzpR+eWgAoyXVhZFw/Pk/et6nlRBcyki
c2FW3ZItBbx3MpVNTlBD58oPGUmTR0MatKxQQ9WAMOr6Mwv7MQBLZEUBc28TR5tcd9oTNB8dMkD3
z249TNw0i3o9jnRYjjdnmtAA6jfdMzvDimik5obfiFtli44y6kRXGwuBsBVIqhhMFZbXD/KkcGIk
hUkpZaXyPUrHiOQv1cdx1nusWZOPYFdVa5Z6cc3OvgY9IEz6/6ZirSI+q9h9jd6c4u7zEFwTb5nC
2q7pf2ZzVQOYPBksi8/jMzlgWN20/61uanxXOAY/v//abDzMsC+2Ls9TZOZTLY0PEgFBaYFbDfgI
CacY6SOcE+mYZj68gvE/5dpgaCqudArdOqNve1r7nM+xw3Of4wGhUZ65xEJJqKvCD1kUUhLIDYTj
zkYpICNfCNzP/T+l0NkAW7NL2JVW/MQSPRBpMfh/jH5MgbfZz2PPQV5ErZo1jdlFekvbmGASun8p
kUOamy//lbvUk40ZF70fqkAhCPZIFdZkTABzL2bfCR19MHzCFw7l37HD8PuhuxhHOo8ey8g/vPlB
bn1n4NqP+S6zp2KeHoVaKND/EFnfjjv5bpIXjp54fhkFkItto2MTB8fEi9MRJl2FbcfhpHl+B4wY
mIZ1mjpDXsP9Ubav/KUCRkW4B2FFOpVnJbMRLrw8zjqlDu+tQ2KA6TaZyGXBpoAl4w6AjxAhXTim
J5YtTGcHflD/e9sm00tICONAN8mCCfHO0DqunmcHA8/EqCPx5fTMZpgAM86hKZhqZKEBKWESPqYC
b5MaWmltbdLoyH1hH6ZNqCUn9Iv+1Oj1u/V+cUc/y4q6L+90q3q0iFKl4oWwZy1W7UawJV7y3Qvf
T1i4Fb900lnRT1m1M54jlN6YB7t6flTeLbotapY91CbUxRQXk13vCwqCJPvPfsyjpv+VkwsJMU4y
SxoZY3RzboYyH3khpe4KbiwWRj2BxWW8HKebnKhziC/4PM0n2BPZzu7C9ktBix3JOX1W7wwPv/tx
2XuzqwabdI5Hwxxj706NVmWlCw1MzLRr8Ugs7keofMJaASrnMyr7rT8oekhq7EqEIez4lP9hqQik
WhGNNBcmTrPBmw0vDke6xgQQSJGOnIaN1wLeKrq0zsK73/Aca/kErKDilFU2xQXWpaztg+zi6RvM
16+qIig6AQUPywEdoCUebaY+yXJtvdlaZoXsKUk8St+vxgAp2MVf5Bl/1ckzLGGCXufXOIB+OkhD
h+lBo7PF8vqZNP+88xns/GlPUMxxX8BLjvFSytH4XFsMLruR+7NfdntBEUDPmFABRR6LrRtfVRDy
2HvBQs948QyCcQ9NObFSCXOyD/rQfPm50cZUETXX1YiJRkSJnbrMpMJXZxTYhzrgwID2YG5cVXo8
YO3JtK7e86mUMhLssT1b+7/v80eaDu2Exh2Fg7JQtdMQrcMwFf34JTYNQvVdrp3vQrqQXgESaA2j
fg8w1PM2RpZ6BSsj0ZeA+oyrPL4E3MPw81l3qkLF3jAxlvZqxnnQS5DGovAEIR3cfE4MLXTP5XT2
gXdsaUhnVA5qLF9X7YATJcx5ovkzGk56yZEnvQHEOIFKzqy0RbAoPT+FUqiY48biZgbgRqeDOOZW
iVdbBK7pZYeGfEYa0HfbiwyKmrQCcx09ePgHhAHXXYZV/CLMmqbxoOneGyaNiIHc2AG0D0yWm0C4
42ICkZMYUYPVb3CriebUVQEP33IpQZaE1ifZtpVvs9rxFfPXWxf+siG95O8hNv+LwCDiLPoUA3WU
YbW9K6vKNvDS7trgdCPsPhihkxwrF0+w7KuZ14hx6FsaZilb/+LLpXL0Om0ceIV2aQKyV6SUgFS7
96gjZTXuBnyN0ysl6M7cfIJJg/breHe4q35OiyJ3aLpmbuBfM6WirfDQWtaf+t3sQq3aKNBEybxo
BjifPsuiQedMvVG1h5fsibw6yfAU3/FqBYvJLripadcKP41WbM6b86z21L6JyB/b8SqlDCcuviHE
H4fSYqiRRannYYDxGLudegV9g76ySfKa5grdTeO19Hn49ruVCf9AGxSM4zeTVTEWW8Hxe/yPFzIw
X5aMkA8ZN+Esn+MJDgQ0zySGfN/zmjwcpAPKL2omEGaeC7WobKop8V8SnuudRjW0MBVgH63i3m/z
Q4FY31eoRwBuywvz6kms4A/95dkkb0D5od4BnxCN3B+NiusSC8ej0beud8QjaDaUlOTzicyHTc/8
/bkaorZTPWhAuVsZKnQGlOr2NhKE/OqSxSQUqmMP6asrwHzR4cut6VZ9PygDcjACAnK2q12DFQ/V
h7hqXJimrdZkeNZqqXdROIyYgTjku2UK1wrCXDZeug7LhFmxaLRpUMUuguTstc0iA+eJhXejJw7H
DqzX19HQmNpa/1BRXcI89filvwgC6Uoy23/U1WWbyUkrKTQ3C/gmSlKug4DH1KeolbaLMiO6uMbQ
grBWgbRbC0UndCHuIRPTabQFA2VygY6QTmqETgIyUdEH3zC+3QNfCGBJ1AD8ou5kusvZ96/VJUST
ZqIBjt54qpimhYQzHBNZTfT3OvvU6Gda+MF4xVZ80JpvxLKxVVQeX+8+nDIcFc3w6/NcOjPJ2VU0
B5Y8PUZjGqKLPVtFVumEOy3P/tNRMIfdXyEgPTsA+6/zavr9pf/7s48dXvZdF6oKNQHcv5IlMip1
4npuiK6THWa3PaG2quy5XUKGWx2pofWtei4SNq6xTp0nZlo8ex7dOmfjuYe1z/FDojW26Zhr4w2J
pTGcYaFuebv6d+pQeLb0DvpxAWO4zOsvChlIfa3e61KyfmQ6qNJ3z+VnpaZc14Wh42AnwVuPFIDa
dU4z8iQmsLFnrqefAQVShFHQjp60eurZj1x2EflBbma/EOCM3dKMbYLi8PZhT7qCgdZcGdvG31N2
sMk99vbHV4zXOBgTGrMBE5Jd42WcYv0qAZh7cR+5e7f4Wcd1q0Inl5VhkRj3+AiYUQ2iHceRgcld
/tgcyQNx5O5TUd5KJpj+BYCzgeGzZvXp9PuX8eo63rbetKgTx3KrN9Hc7qCgUk9q9/FaZzm5Yfdx
GhIfHFf7Vdmz3XNTw9jK5V+2vRv7ukT9Ctx9/a0wpcf7T0op+atbFB7V4Tb8ClHmvewSlN1Ahw0x
w7mFdiz7+WTd06f4Zu9ShT47jm5EUsJZgS51pqtZpo0u9ASf82UXaQ2FIY6ufin28dH0vuq3pTG8
I/zxgSuY4rXuqXqmIoFNmNw5ZLSk5TDizgrwrmzsH5e+yteDMH8MgBvgoazg5wijUVmBHGxNFxyx
nShCGX240ba98PmbymaIO1yLOh+W+2EEy4Y80KGzm14o/SXK4imHSj/cCgb7AvhGrep81jVoKeU/
PdXHtq6FP+Om2RWbsmlNEDnxH28rAoLWSDAo30z22xC+Xp3NTfIbJ9TZVgSG90m35tGIw5mOfUdt
vmjreIkYX45XSX22ko+pR1sr3pLZopA5E8pYCZ7dg9x96X8AikKnlcA4MfJRlpT9CfxfRDfFGvwR
QYMMSxIDdN4mYTfkSOEF0StUiKOFZyKLVTLdXjXgr+RIEUfKFKlsXjCTcN/bezWpL7WMrQk9W4Tg
kuMCMhm0//jleYcMPa04Mrlvrg8lvZeO1ucrv7x+mWwFU7xA9MIBMehVDv2b3EjTLd3InZcB6fW7
azjYc7a0bdNCmJ09Pv/egJuQkNtGw4RSTBUtTnvgtK3jcplmeOf8Tgw6cuHx1vymujKvbRbAPfqG
FzmT7kK7wjEosTcUj0kjJFjfhVU+w7mbWtAs9G70sq5x2hHA5K013Hc83G0/tgFoBM0cfAQ7pU7X
y1MfJvkiGIBy7g2so6J3uw+XXVA9O4fPPQbtPH9h1SgN0D7y2o/XeWncGeTEHPBj8H7c8GgB8fgl
YrvdCPmjRy+174TpiYrWPBuqW8DgfAibNkJ96bDG+WZmNNihofS4ovgyljLlcj8YLT7UqYFr+1sX
Jq4HVeHG3wdT0NkGuA6o7fpsVznBBVwxCmzTBMc01/vVVVHVcUKhiob76ZFsDpxIwzeAIpBdUdi0
ctarufiqerHgFO2E7QFVaIOEBqJuycQ4zENmcLA947zWZgvkSILMunzrseZnBkaoQ4/CyGnRrx22
V1rovijfXz2Skm0XPbqGpKD7ZiBgdi//BuFeIjbOgbMd9uJhBMNhxjntd8GNJCX7aMAFVvS5YF/7
0GUhkjVPPbbQcpVmQ7F1XAx/2OsnMDhpt/T1VIc1CbNPell1ov1BZB6MvvhlomHOEOB/tYFHtvP4
FUAJU+R90hjCu1j1+omhLFEK/5V9sj5zbp8f11iBsOnrJotro4GJeEIQ8A3hFxy8qNyJyB8wBh91
GbTa0gAPgnxKz2msLSkcnzQJs7c9XFiaP9+E4l/fH+Y9Jr6M9SURNHP4Ojw2rJs0If5aA/haT8c3
ab8JIluAVf8qJKX6qhJRln3DjQnfCFcE6BfRLKI9BFeuIPdslmGncMxxHqVpRH1gdUgyiJeafP7j
izdENKLZSegB2NZRptL6C8jBcrlw3sG2sInzzxbOLWfAdkaKaQ1IzajBjeqJwIVRBFBXPZa1Cf+j
MQoZoABrciy5E24SeqqXUaiN0AC6MI2QSVkp8PHJHGhfiEf3VxiMO+tYDJlC+A6RpVIHzYPj38Za
F7VSoqnsr/03D6d86zYSsSoOdxt1B3+43bw2ZzWihKKpqcAvCv+YCR0M5DiECLcF9RpccJ4VxCNr
K/1Rx784qedaa+Qt+F6oqW9+nt9I3CgzSumm8AW1DZLLKRGXlG9OXHXiUeZL/5mLSvxEKKyidk1F
IRWLN8lXg3uReVik5SxC/y7vzgNbg7r89Pq0KElrQDhQgzVT3Sxtc+KtxqZ1P39vAX/w9UGg9qNl
xtyIp9V4ihoBxxgtvrQhpPIf8dqdwfqqCYTIsP3NveTzoW6i9OHfFAuGm5WQ9SX5y+7rUOHdX5ia
ttkwYJCZGtwHBQ2do2ysMBbi9G0goCMXJswsvRHfWhxlJPloOPdIEh+/zVamzyHW3D471mBlsqbH
uZHKL18M7knkdtYvfG6cZHPglPp3THZo7TQbn84ixtoxkZl03OKcOo59H3xfpI1XkYd+S23SlUw3
q7CC9zzeMwqGjGkKRvNTG1+GA+t2PiJ59LsnkFKuJ5TpPJfNuVgzkz4igcIiYEO2Dj3c49RfIp8g
2kf5EfxH9zHj50Z3hxw1RFeiq303Xcbnw4+SlUA37wbf6e/B1FrmB1QQpLtDh5BZBnmgIbTctJ3J
Lq3+i7LmwsV/unoS/O4CdyKvyLpwVjpQyXKQaQStsyA94XSubn6J8VygJGfNCMfDWI/m3zHRimcp
TCgaJNyIkbgWrj9gaZL1C2cCum1RxyotbbQ8n4AlK2zs1/B5+HDCtwTRjP1HMvGBwaq0HVVhUrVo
hECO4c4H8zh0nIW7fzj59XVD5p1Y+fLHbMCto1KshSspippTEWJsiencs1PHl1svoCGdHtFr658b
N3JCGsAqrzefrUQoRcsmJVbCk3xyRsg1D5/RqdAohS1OlTrugJCNvQJ/GbZYvnPli0QK946pU5IT
rhmt5rAJDOIZ/nns99lAzR67NcKU2OsqiLrbfGVERhHrOXupuDILMdNKKBSpka5jDq9Fkgs+wY0a
UgSP9CQ8b+aNBQaRQHnQmxmPAtLTJpRil4K76jB5RAwNN4vGxdDlfkdrPFP6FiL3iZ44PFOcEEU5
rYecqwegtaP9El5Wo3Ui2NWtRxwQPm258YU4beLOu1vHVleX8QXkuDy4QcW3x8UBGmjmmpk2K5Ny
ev9YvO8dhPUq+JdiwyUDdbJVb5sAnlB+2I7i6GapDURDSC/0DOUAROACwWt3a8Bahj+36rJY5D8c
ddUGsQ3+eYNoSV88X2Erg4hNVGgNN9soQFXEVTx2POP5ax5ocKn1eMpJ3lvEQDSHulOK/D7K1KZj
MB5awmaMZuT9HcuWrwWBgSR6XvCqfwpn6I8N1qEzxapId6/yLmDuTN0GK1swbQgZNc5mIrlc+C6e
2TwyhmnXHyQow6v7Bbd4/HI+pfEuLkCDso0eA0PDs6db+l3pG8fAUVLbGUGlip4TlqOOTsDo6isR
NEDNDXR8lj5oo4r47HYg5c+F9ndReGKn9TozJJklibXEjmRX4BVeU5msLefKOKuf6LToLKC7a1FY
6IAoIJksVUFwqJuB87ZMsrCXNSFpHpr+KjyP83Jq6D/K7iSpdq+axdO7t4ViV5FEe7Pavbb8UlJM
NH+Ak6w3wz3kA6+/68cW9Rf04baFsst7bf84Il7+Bz88GbFtsEAG8rrhwQlIQKOIoH3KCC7VCv/c
pYC6A3Ml5C67Vwg1ks/Nf/H03+1UjexpfUbXS9k4YKdNmLg2kk4v2gwMx/wR0F+qZBhBu817Aa2G
IHTrVW46fyIWR/SVLlN30LvdSloOo4FOt1ZTOOP5clu+QTncKiuOxX1z5Km7tFfgYViXBUYENBG4
v9mLizpmtT4i8z2mvmzrDx1lbExo566SpvxVRMZGGpThsXQMQE9XDqz4Udh7bwO69rcxlCrFBPlD
Hm+HZNHTYnCsWNSHcEvkF3vUoVsa+PoFuAv1y9TFdShUg+Z/2dud53+eouV4rIInQo8Upwifwczo
kauRn+xwk/FEpGmcdKkqICqXFR+UGhHO7qww9cjSTdwR9bblOJHjf/RlxuAHHSabnI8gshiq53wy
pvFmXdmEPzWojOHARQ3WCGYq7VRdH2HOysfS3h0vXJwL7lfX1ebfKthmbPV/KSUEnVTLPZlSytqh
58LFg0eIItXQ70ihMWAqfToxb+G34CPV2ZXVofD5aim3K2hGh9QVGTGKT/kgKYG3DfVSWZDPs1n7
WZRo0JTOAuXNP1uys3qAcfyYIqXf6i+sNzkQZ5fAaW+A0DBpB7CxFN5hRE+XX3vd2Q/CYGQixsV/
a8j8MI/YFjO4PClanXfeOQw8cGI2umvVS+Qa4T/9VYp3+BQogn0tFYI3uapXcafboN2FRKn9wsgk
urzH3gDbDki6a2HNG+Hb09gYHBKpxLSNneGXlKmr5r5EIgReIpxk34m1r1TRaGz4oCQpfZR0qq7+
rluSj0gCtt5cEPPpF67w8/Z8uCeWwpfyWB25HDoo5kUg5qKe4czvtz02hDhMgwSKo/QEqy2ryCKb
z5z+jTi8aUQGwjH1LJtS/9s6PwxyKGIAp+E0R3BteuFu6kItIeVN9DWmSFCLaaHVJ7XsbXqbArAF
PFgHuQm8MovpkBFRPNotr/HjE3yGufBLx3c6U0TJbkzW3OlS+OrPRyj/4eaSjLyFI+gU+KyQGqbh
8yOL/lN2TWL5fe6Kg43sL0uDJ0pUCkBzfmQk2TQ0HVJHIXjsu3N5yIUJ0ZpEg/Iq7+VZbBFZLO0q
E92Op0Yl9KCaZnaNrDCOIV/oRvAIRYX0F8L45g/l3djNxboTGTARS/ahcSzse2g9g7fbJmeEaoNV
Y2uqBNqKLX0XSk2L00ELc7uhuKDX77uAx/nOEcIGtfXkOZzsquRCWikpKDcEKlP903lV3HPKh0sO
TZJwIAcq+wC1dyDMA8rrSS2PsI+Z/VEwAAvpB4iyFqqNiw48i264JQgWSpag2yl2y+izSeI0Ixe+
7paKJx46umRyq9YlUabDpKUEgQuUEJ7Z9ZUhfecOTiWNnGsrCJ9uLnuMVL3qXc7p2zfP7wE3SEDH
h7CQpU5aaDCJVIY0axNuirhJEK6Kf03SjVotZEbjVRqOaVIao9SbGTfK6CqT6KikyrGdym8wvxfq
LRH2at4dvPpceS8PU9g8OolK4ayguyHuJjrbM7MUFC3LhS2DsQHpJfsyD4pk208DelINcPABc4WU
79ySWbLMinCApSQTYeTzEYhTYQYOqDUumV0Lw7u7zllHtMArUDeJ7aLkZiHvj3J5LM8wNXjkD22v
HCUHzftq15TfKQuFRCsFXv6k1LjCb8MXdcnxGlMOrIyA2DG0cCs95pxsyg7iVszIEc6IryKLirLG
Tr8r8S4fAzkH6MU+pP3CA/ameNTgotQdYPdDPXdzf7f5917wJBDgPT6fyxLSIpxeETJf89CiGQI5
RMWxgrVLg0qhyv+uRdP7Fnohus741JyMF+fGM+OUCb69qb+qWS2fwZc7KCwDzmgRYUdKtiscGRT7
8cxW50QKcQpv3AInoWzlGbWI3jqIAe5qcSjT3R0P8295poekECNAQKlyUtH/cl2W6I4gvpFb3ifZ
sQMsH/k6aMYWbpKDnx1hoyikW+pNqViCCwtlQ8WMwWr/fka5d3xXGEvVc7vcUIV4Zz/iyHPiQRUJ
d6m7/QpM2OpXAa7wovQw9/rVO/mKLMPrWE5r4wozWwqL+kPiDigk+BNHaQwqWoOyCbZq8ZhkGcpx
bgMPFZb6g2UHCbDjfBiQbeyF1KJEFrHjlZVKUSe5ElkjMszu8vFUwptnfViSNOKNW3Fe7s5gIXZu
uErlDvSGaq0za+Db2s8Fw9LBc4+iZDmOr26cfM4umTdiB5bl1EGsN1mdA1eylg49K8os59+H5+kl
VwMLQUxleRYJAc4IxUkaNMoDPsrPmxgckeukJwlTK48vCEFGKcsQKrJ4xpjcXsBXABmgrj+DQ9FQ
0ugOP23ZzwR/Px99L3GL6OybthI/GjWENZn9ZLHX8EGxJHDmcapU5C0YvdoDGZkXGWzz51abgUZz
1nB8UlFzBBgbQ5psdV7MkUo6Et8SzgkZxrR4XjJRVvBdS9KHL8D244x9+gxhh3cGYJHxkPE2oAEu
bIjJn7u+3mnAGXZ4PBJSNYWWrS5tU/NWNYuk4ofZ+nkWgXjbYOJihFdnMzL8JHUCQyzmiBG4wVdO
V5bWArzB9iqfmeA9w8tr51RdlOvmm1msuUbIiVWbvNGFvm1Xm3EMGtpx5ZyaQsVL0RgPH9r0qIAM
FmuEyEtDT+XX0kkxNu9AvrSLsbKGq7xaREsu71+4Vz0aXAKKEzEa90WWGHjfIy1qvnxafs5c1bwH
saFecvZvuHgu//OFHS2EoydR8+FEeKMkZeNP58Y6HSCmuYmvHWrc8A2kKp40c9jAWiScEsQeFzdB
yw6nIuYJ8D4NQdiM/xK3ONy9dVs/BgwkimYYpMBotdcfJvltPIrO7f2hJqm+64mjX2YeYx2/mG4Y
u1C0C9CPdwpDFCFQhY8g2EIYtH6Cv2vbBeMf9kJ6/5JX0WhbEJaZeRQTc+u8x9yQcBMyEH01TLSc
DJ+6TNs+qgzEqN5pXntwxJYfP3J9kO1QbPFnGVNvAmspkxdpqQBW1l6rSt5PTAsxR19elG73XFEy
r8Z/FpW0hN1/6CUBTLpQp2Mybv4ICEwRfwue8WojYpHxUyb/+X8VjJjScFMHJFjb6WJCgvmFJNZS
f/QHQML8pCIqOSWiOqN9YR4CEytBVqqp5ocHN8J1g0LO6JD1NjkQ1eJWEuynMPdzRlo5mdPrO6Ie
/2iBUEBL1CRDJ48LRCuTzljKYapgokMHZa5A2c0EFvE/mb/qdYhpW8YqTEgV/ZPzWIfCrOcNEt39
AfkBVd8AI2HrEKVJMz9YF9QnlB1r/QXSLtwbLPGqnt4n77+2W5bkteFNEdHBq4pAbOVvshMvPDao
18HwvXbu6P6xZTOvFZ0Rw3qRd5O5d7lklUVzFr+4suFuQcOaQF3IoT4pq00cAwiewf0dTK9bz/93
PDvhrKsrTANMKZYAK05mXpKRGNw3yUBh5OJDNriwHk9dl5PihNHL2o0W1WIgRXJ2SrcLlazf2lO9
rcoOoRbHtx5ESZow0pNxHLbwrq/sIctbotKy/PT8cKGk9g/b2tMc5uEFc/PV5z3Y25+VpC2DA08o
DmqKdBNrVUvmF25valgUDmH80Vt/ARl/jzuxVfwEyAjk1oOWjN8foL1KfSYKwmng5ZwSfbdzUj3X
3Neoon+gTXnoUhjwUUP+6IrL+yBD5z9yQKHaHPQam/8zLrg8iSzfBfsKzPedEd/EqPbDnNyX4nPF
y44QqKViEdtRGlLHfBWCYB0QsnTnBAgn1c8x20FR6oZPTdvrtPZ99+AE3zRJAxc/XTFi8S1CYEhO
B+mDX/0Ud+FlX812ay5CBpvniTInKUourkX6A2HrYBHPKh6LOEqIfBIP6CLxMNOYBVGjUSDQXP5K
o78LfHk9Mo4FJmT130tA9mm0OXyrUTGE/ZKe3WEO8x+cMpK5D5IoUAS+lP2yhXhcjKn8C2NzdL8j
6Waf10uy0jq83ivXy89PvSmzna7hqvJdWdMOWhZqQlaqmgUOfIql60eUJdC3kBlYbTlslThToG+y
mDj52aN7xoZ08NZHnFk7gcUU+D4c5lU7mD0X5a/Us3aVdWXJpI6EysDZsr9gl6feSw5MRBRnxCLE
zPwmZ4HnIng6YMjijSLLoG67bHsEjLLiubukHydFbHvzGLlhCvZCj4WbPahQAZBu2QswrhEoenrs
D7DBs/Kbiojl87ErUJdmPNo72wWLsCx+jJNW/MsLGmQz7QY3tkct+kRIK7Z/RHZBbd0CQp4S8Nrh
LwpR7duFBCEmj4DnuygWCd7MA7Mw+eUfHc8ps6Uy0zRReuV/+4pmSRDm7ZPbEwHMeU5YlQdG+mzz
JlMT6lSFKcUs2EL+gvSLPmKZZlez/YYRmT0vKC57Y45Jo4+aRzDtltvmAIuYhb19wn4aOktG1j7W
+BUnkj57PqYwFps0dFDNIs5lmpkIzKin+WLZR+gWW50wHDPyx+ZSGNgo3WWZ1G1EB8aYF6sJ0cqk
CWDe6YY1W+nLEXGI6PfdmdMouaYEeOeQDcnAKHkCQedliEo/aFCI4Sf7wFaUw38yL/Z+R29m1Wsy
DdTeie1M0KMuZcjLPxH2LNdnUU+eyJLf7dlumbh8JIGkEfNB5W2VTL4+2EvQ0/TBqn5Ocj+kSz/k
NSwWEFmFQzvx34lf+tZ4v2oarrWXX96oM9TgmubpR4QN4fTUd2MsERTpYR1QLcnB5fNzfEWahC82
nAEzGacaxpSyqXMXW9w6wjMIH9uf1JOFMAAySgBKRwyWtI7084rVoQpMpHHl/Cu46bJyEY/eMQQR
adr8KrMEtr+gkWkq8uhBTSzirocxiIoZz5Cr6+pOr8lgzm7hx9T+X8ogSjDDetuLCVz3f/OkP3LU
xdAsSQ1Qr41OAclXZzbW3HJTHhkGeMrK0BkrTIHcJ8Ys3Cdugy46NavXEMrG0ma599WZRwzdWxq9
xSRiRru/4bmJ08q9Flpt2XsrAnXeNgqdooyb4n0dr9YEEMZF4RfsMvXNvNfWNigH8NMxebMCRZTz
KZlyiUauCmyI1UQ8dPWOvifJ5XG5KjcOWWTKL8u58Zj1/S0ApTQV9oP+WnOXgol0g3WbYCEJEZsI
rCm7RBa8LVWH86PLx9KCuGDz4i2TdJN0ywMDi69eF8Wz1ZTuguGFCBfhgq4cOxJRPPAUvMRmD/P4
UVjLJtEflki+c4MfnEAA74G7ysCzEJQX4vkGrxz5MGiqMUZssW8X9LWjIvLE+awglsyH38yA6rKW
iDYg5B0NbImsYQGgRoLKFtlesROw/CvIu0laymXiyxGIAfmm1LAWrP5cDepSzUxbz2MSpejJYn9X
0H4GO1k1M9qPjpofIuWrwv+FEmlcRWkeJlcY1eF8+d5Qp27dFiRe9MjDicT05dmF79VQE2X4K8bD
lB9ZRm3Brr3vaNqwqpUSWjVRjYF/iy2/Mr2dPWe4Vgi9WDG6G7rWbpORCZPDqE1lbNm8EiKz0lEt
dvYFQU47ti921tTwaXVeU4LKsmD/gMGBPF7Y4pUGEQzkPZrBH/Oto0Mv08iC6HckCcJX+1u4c0G2
1d6g7hc3CrIMhnMf0AAir6Q/Mepy3MMZSU68khSmyz5TtwGJ4x+u5cnKns+voa5QtY2qYvk6NUbu
6gzuynQ6ZIgINGROkwSMmdTd275M5qm6fE0dqvSAmvi2iktZjnjqykaUpfspqADY4q/pubfspzR2
eoNp1ikE9fxTwZIcxSKToCAT/CwwQH9ZJCxsyl4R1cy/QV1hBI/uh+HNOoQfnH3w44krpYgZPRF0
kfZswQgtr7wUdM+BCv93jIY1uOON9TOuvw5hVcKRFVzgxh7n3gdMtDOECNEGdnsAoqqHt3q+kiwy
0mUXGuBzF74OTXtCnm1ycjPFiSURjzsQiPWKl4kvAhULAIhIC7zFNsINUl86/vHZCvgaMRouFrgG
5kdPpeU4o2LM2Ozksx8y1B7ELXF4RO7xX5G7wn5rENoproRGbdAKmAvNEvhJ287qYxkEstaKN5Vh
v6tR+g0LHfLoWyoZuDbfN8YsQQ+GcEPdPiJehfRC6jty9zey/R1/en3BsGrnE74ITIcZ+h5A/9Mb
/kqbmkZJtOs6c6jCx+lcazOlTxm5PeIHDenqB27IM/P3lndlT545Q+oewPUfReuNvee1QWPvHM/x
kV4g82C8ObKup9LlTe4YGghz8W0DBvxHAu1DxoOiO2J3aP8EI0hmwENnXsJRjd82hSFjQYPyTTlb
uCcFBj7Frqk5XOEq479gO4FSjh/ve+/WMSE7LlePG3ixJ+aBejJs+EnrZfi/dC3yw71ilsZZJDzR
4e/yGV9kUv+BU2N+FpHIcCVyf6YDSxqzeVEcn6tw8M6mhezv2rMWmwOYNm9RzIlREOc4cco8VecP
7CziL6y54AQZwodyYf9FQ85nADMoM97XrteyNQnoe0ntdu4oyzNs5+XqfFbeujotlB6NByDCTYla
el8cKFTfckSLi9aWCM6o4Qe7qR4A9VIb9ElpJbpSArhwSITnOmTYU+9DeudtR2TCH0vPcWWIpThh
1pcOEi8VfcoLdGu87+AceEC8VKtv9x8HhU9nTRmBEhGvS+0MizU2RjnPA9jRGmKJvA4HkugibJm+
acP2X6MHDMXgi0FGohZjuRmmbk1FVIFcHmM0nyM+bfmh0JIPCQ8M80UgtkT7eOkgS+8Xd13IVs8d
Jk89qbD0XNARDR2NZR1ycHnRBUB/gXmddQjZml82D7E1njIz3hYw6PzLZwW0Z5yv6GHKWil5L68b
pp9/Ss6Cg8VHDTIxQt74ztHkosg1xXQbe625X1m+bcb1kStV6vi8sUAtBl7PzLriM56frdf8s0WP
JqjsUi3Q8ftwCU+ZF2gStTk23lQ7QGOaAqFAwR3YrLsQYyeDXTrQDF6tiom7OA/urRtbkCy/k60X
aXdqtgmc/XPBEIlogMwJuyxH6bMdL4JR0CLUe2niAtMAJPntZM+8t/NYP8YlTF0WwTsOJFK66B5M
sXGkkGlZRve62BY173c7lObl03jCamSRUk9xz0k2k5y6Ow3lKPsYssNnJtM2t0I3wZow+jNhB0Mz
W5rhP9WHqUpd2FeVHFw+n1f98f/vpUjPFkwNKfaGG51q/Q7qGzz5eC1RiEDxRYFl08PpBnNg3ybd
fkmrfuxBZktosuNs6gT4+eoVLNhLdTfpRJhSJGM62DBqPAd/HMY2Alh4sBCTbcFRuoM+KDbBZ09F
5S1EsUv48oVp4fR3yMZpAmikWpwGQ859DTE9QplYHfunPSiM34qhBcJt1dVnPUsafjwxhfrkS5mJ
bOv9Kp+w3yVhv0mw21+2tu8cQWGaoP6lHR3rr7ft6KpbMByAONPxs0afdvptRnSJW15zIZ0Aq4h3
lEO6IHdFkbohmK9XvDpibTzfZw8fNSW1zNJysJHiN6xYfHBhru0A0NQvnqTg3rRTvRWeZuKuX23m
MO4IM6KTBy7vFM46YSwtb3RE6CgjlYALKteECncLZfFl4S55IAVM3t+tX1WDHF3s2/qnAWelf0wC
1O0ygwOo5ktlRnqeFKce5c3p+MJblHDYv/KfuYqXeZBvs0TzdX7Uuy2vRpI6YjWAffYJ/ch+NjdX
6MipJ6c/QG1umCpYsk4x6v2dIuNtWQO2P6HFJujbMS2x+jaOsHgsNTRx5H9vDqAf63EYmSsT7C0H
+MKAE6yIoRBoDMtxuMrjVNUBmJphPro4oo1dWT/7duLor9T0qg2JF3fHCbxhg44FiEk/aj53IIE5
f0ZLd7lu+3xwiZlT4i2kBmiC4j8Rz5xrmkq2stbrcvqWMNTzaxuTFJtNh5HRyaJ01/AnHFz+KUeR
gLf6BF/pNeBZyiKGHuZ/i7/RcuKM3Z2+n1pofoq3f6eC4rTDtp1bDNR5yXPdcu/y5p4yfUqqYILn
r9zvEk4s+KrqseE+7uz7LXOANsZMWIdUqxKBZOlLm7G3tPa+wMbZMWFvl2Zypml+oaFJzVff6rhK
Qn140XbVDhRXVRpTfmjcsW/38tdhbag3tEA/gdF+Pgb40vowEZk1y8pCVwaU3RILsdYqfCPE6PIh
tSs5gjg6z1mxiplUcKmXjWglnHd9bUyIVF5mokG3s45fZgqHU5/O9msSsszSf5s0pWCTCWoPJq9/
rci4YqBRcZqug+N7CbVhidk2Xz/7BBnpNFJLW6ZYFekUmh6Wh/LFHeoXb0FCgG9NPd+/G/KR1Bok
J8/h5F6pUT9/gsBcvpaoPBhm5GRXV1UNLR39O4Is7N29Tpf5xh5IzqpakJbZMLWySpYyl+e4toQT
Nm98cqzKBLhJhS0M0UlaKpRidKRvP9AhCes8EzKF59DpzEy3yhtdL7Y6iv0KhQtPbYsXAtaTSAf8
CkkjJgM3iSXKbIgeOGK3FwH4BWsrsZeVs+FLynF1r0Mzz+8dwrYUs7EfVtiIMT/2KwLn+IA7DlBw
lO0HPeVtEegpgh7Sv0dIUBqetPtYTfnFdDNLZW0IdDtG0GzrTXzes8iEKIkqkGiQCxNOYAGEAyj9
vqEI1JQ1TM/d3MmJc8I8Ntz4e50f8u2YTSAFdblBYvAYWVAjTb5BXLOCdqr6sbjMFxcSm3qSFYdi
mZZvrWALQInLztIX5nU7jHb66nxKGWueVewXXYjKnGDSPnPGpKvS5KcLoMsfjiR6XmblD/p6FdCA
8jLVAs/OYtdBCri/ShsfwJFoKGcRpBz8q9bkpLXWSERbKr4l5jkCzfN87IgAG1ywKtqg9P9+5XMD
6RSk9pPD9PJZVMoAE14WWG1xcTHdYSI16WJ6TSljUssGGJJZ5tiu6w2mtmMK6M8jWWdlmdV0LTVH
BD7mvEiWKn22kwVj1wIw6MypzER/thsn15GJrAB4A2Ple/OSkLdQQyWkX2QPd4y54JYe5YsVULC1
bnzLRMctdLHMRtdY8YNswR5mGregp4wiZPLZdz8WftSgQxnnDIHRzE5/rmW1OTLyDWZxHHOF7NSX
cY+aSiuUgBQ0NbXU7+7YqvPJpGLZ2vRwXz7Ume6FqioY8cDOccJL01HSYEsbvg+HkfYXG+arUgmE
N+spdgt1dRCILhaHI/7hLG5u3XJHkF15B2Zb+ntnXNcN+98YW54L74h0PdjY9Kps7y7ucfTYGKew
vykuc2QezfCU324Rad0LwHA9SY5Jh/BHjIgWZ4j8NOco8Qg/vy3l3f9dF6J9DG/O1H05ewjBSuck
TLcBPxjOZ3jfXxpcc6DAdisIsm48JQI/oEaRQI6nwcizw3yLTFMQExe6Ck4aMol+aWSEdlhj9WjF
4xXEdZmfGL7jKQbW8XJx12eFWi3opaCwuIP2FHYg7b4AT6FvtzqZMy0vFcMIxNh1onvL4zgpk7Ud
emRgxOtP0ipHQzsMuPupXtBfvNwpd628/YavOZFhwck7IgJi0tQs0VYkOaY1xzrX+OArl3FQXMLZ
GqEP0Qu8Cj/Y7ajlQh/X8Tcu9qNdinCCU02za971+nQtf9XB8aiWMssWP469fEniBXLQaRjHbPZI
nVPSF/OU7iJ08SYz3AYsWfeZ506+TfT8xGYS82+U0p3js9dy1Rinuu+HtGMT6eLNPyKLUOD45kP9
74tYG6G0wqn8jrWc8SOgVSQMst8XZdZtG04VJARKVLqyAdaE7x07PdB34O6LDOZ8PuR86Go7Us6E
ofJL//Wpg8nasK3Mv8MRnfsCC3XZeeHiSxRB9DUVV43DDf3nw8/F5LPItyYIjOqihUL+gFdkixV6
UzGCrTxuJhHOJMmnVjMIyzEKgfaF/CPPaJUA9tIGLuyn94wM0lpxhywGtKiU/H7Qr1Aytwf1gtqx
p1SIzFBsEbpTcXtw+1uWFhMo5PEohmfQRVOBiG3JI7Uu1e/7ju7WDUMq6MImwxAkpZ9+U810jHHz
OBV82+x0LhAuyx9fy4fIOv+aEv005/joPaIb75VIbubokFZlbFhcV5uHXoS1QsTVOcHl/W0XEmrk
1vbsiqizV51cse/HqTGv6Z7VoB4moonxGaghdjNh5rwlRpt/htWOW9mAO/nV2GpbgZexT+8OfLgn
PrGyQ4hFvTEBeLqO3PM5cKM37gl5/F/k8qFPVew6qiSLq++903IvG3NvOMBhHDT415Sv5B6jsaXX
ShVofMrevBgr8wI2U4xAfqyOtkWX2Ns0MXTYwPL6iZnvjLB3XyaA59PABFNv+D2upQPFUNIigz/8
80S5sBq6EhjpMNxNALBBDQntr5Sv2otecb5I6GiqmoNeStd+plsprzsD/fxZTcKb4hAXZLL/yydw
bgwcSJ+uxF5o/Wmhv/W6J61weMNx5XJPgWl/1t1Kp3rKTOxIT3eKlRRmPF/1+l4bcqqw4XUwq95K
/lBwyIeFy9mg+FBtFhkoYM9QaRBO/cktRW01iuCB4UYc0GzspnH+52KYy8CR/2LDgMvX3DT7AYBJ
U2bmvmPwA6pa4xFjc0iFpQ58f9J17z1k8Waf3JDVvFHDAfZeEB3dyOUpFQ3lnnEzP+aPynFVwguw
ipGOIWvC13uak1OLwDV+kAL59ygMOPJIVc1NmU4BspnjrqfqsU/no4R5gphvJelmRYDSBCSpX+IE
5NEZOchPa1cg9TKIUVfqtuLgPkPrXBBwa2ApHbQBKpMpW2j0Qo07+PhwnIsywLQo/FzJb5IQBj2G
AepQHBxknQYymSG9uLOJNMMO9zcatWMxGaa19acsZxxysmjelgROeDkhAXlvfyiR+LF0dKdbip8x
wViz68nvWgZXKebTTXG6UhhOYrtBLkbzyfS5v/Ham1/Ea6D9TumfQM3K6mlClaruJF+K/4CJ7YYX
JdW30Wh4DxDSL6mCyJmkgHwXX3kpsNl4RwT1TwKQLBYpwOs0kKAhtUEhQ7xYbMSWakr3ukJ+w83h
VbRYI+CjRNlGMsnggKpIhs5zi0eMQ2yJGsiWJncoAgdqW7VBy3NMb3WMfN85aZ77FoFCe0cf+73e
jUolk6qSU9fHXhs92rEKrGJhYVqT9bM5eYHzRxitrlDJg6w4QjfzWHHoST/uyAXrHpXhzx8DNYpj
HzDbcl6zXfvTajICU7YMEcrTVOZXj+oJrmjmIx6NSZF0EvMDUgPaqYx4oylnnIdKdqyZvOlH7ojc
oNz+nNZ6s8bXekSHovEVUQYWXflHaqVSZyKOAtpVCG8BTMuFNFilfHBuJWig6VXZTe7zSWldW7bL
fMYvnSN0C8H/swAUeLjwXU8fEa/nFQYhey5y2Su0gQwSroZMrr9uDSarkTxXN/3py3Ixnh3GYtYt
/N2ROTaEtw+5l/dJ7xyg3Y80r72MLwYTe5oypUFKm5OvmxnEnfOC/sLd0JWZ17KztbZPFvQR+S3+
o08LGiWmLV6DQHjpbk9iqcgMxvEISQqeXuJBjNz/E7R2YPCPb/dfVlx8tlXBwlvw156ofL7O9xFo
ou/IvBJ12JXNNzDfGsmUNWXj1x0uWYXLqO/PZI9XrXq6eOcocZepXCgvzJzD4jKuZKZJytw4HafD
2zzz57fvXPubgaSPswR2iV/gYcUtvT93Fuu/N3DcOQi3mw0ajVzvk+oxRvzWcnZNxh8P77kUu/fd
JNRmptgbwS25k2LKR6adsvwVO41wVJWNe+mGL+w+I4iZ64mWGLjrSuvivNuBuU9+lOQYTk/STnsu
q7+xzsNLDTsuF/FLwRjRqldr0p7NMiBgpbFgw4hXA9LUqeSagKwE4fSCrT2Fl0boSTuEJRkUzjf5
yE7sVpRqg/WKc31vAG0Xk3I2fWN0zQ0PhAu+xNKbCRFhT+8uoaa7Pl8e68KdjfHUW7vrSyAepIb7
7SAL6FgN3EoZu+SgQkH5vgy1gcJlZGShULlqYXPOKIVFMEiosx53cInJ9xObthMCcYfKELvpFWOf
J9b24wPYggB6Un3xwpu+6GpUZ9V5l9Xi/3sEkTEKdk5oXezfnYfh0jnKGGJwMRL4eBlIBc7GYRow
m+Y0+PQztrLQbBfI456aK3FsJboQFjWtXw7L3trdHlWNjR4rWMGYeLL6BAuD9MSTAdiyWyCMjkz9
h91GkGfUD9CbWNpcjCeyk/0qqBvDa5v67NXBBVTB0ysCaJbJUvCrp5kcmM2pzM+yvK0I+FKFJcoF
EufZ8ovudNDbxAEnLyv8NIADA1fSllwViyCZdnAbSYRCYJ558CKxfkUgUHlCTuTXLaEj3B2WziXV
4/stkzsyi8O8qKX1eabNQPfuxNDHfeHENjcZiUUeGWF1ns8OtgFXkfDBcsK4d29c/IZQSOpwWPgx
Y57QoWN5LCoq0KtNha79py0UQuey7BBGWV3XbsbOAdLLDw0HJIWOJMaY/n433xKS3GA1f6hNgDOx
rRh+8Scx6ds8f+eaR1Qq1jNOIjECvTF8wq+4kWB+B6/JmglCW6LOVqxqsAlDN8xPzh0g05IbHiq8
t826qrNWRr9VBDPuY1EFRo58Lv8b9/3OZwqoEun02iNYqVRMrLj33BVrhrAchOAJxT0Zfxh1H0T0
K+umrcs71iNhHWWco92XA+7j0BQ2dIRk1qtFZtUhTXJjRjjB9lMxuWlfnDt/IDWeacVDgUN0IdLr
ENw/13irwDWNb06d+G+qShtvFjOCbEQLshA2M3Cp33HJ3OgMAhCuiWzVHZR6TQ+X29RDER7Wt2O2
eChJ2sc1c1PTdmpOFTmzBhej/HVHvLjtce9CyoUPluiegT7vv0ysWXlWC1WDU5PSiBxlfYQk7H8N
9omLOI6+Jcppe0xN9OeTMq/VUI3Bk8C8LPwL7+TBUkjMZ+M9Lw5dDVXFfyzaUp7f8wF8EVN82PrV
2UHNfpiFRZkKUW0F1+pwNLN5T/Bpg2qJ4QXDwlalQpjcvEynFPk9Q632w4fHfNJiwQ0FGfnuR/An
SkgCMWDPTEYET4XkifDew6ohaGcauh2sfnd3jgrRExNXIBFcOR7SHZKpCigMZPH/zRsviEpRZgD2
bAtMKXj1qFkr9zJ9qeYuJ8UyGfTJf4o48Uh5A1ecL9P5YJIFnuisNXZo8JLz0BTVTZBOe/HDGLAq
YSx/tfe7MjdQrHzBpUY7qzHri4fq+buQsKMK1Z9opXul0HT73E83IGzTOc4lk1Lbbp4HqYEu6fSt
nDka2IgzcSiALqCIpSPdMM6QCBvdCNB+QZU7dUGaYhyl760o7/2ZR7JBcFOUqbmgqGhF7c0HQmh3
4IzQbBJX+8rM0NJZzvNJrs583IKBP68SD91oHbIHBllBOZO5KaznbEsyulJegXS4p14/K2BUGXS5
IVF6Jmb8HHPFm7rKhkcoDi2V/5rOkQGNTyi2XaYZq5Xb+CU5dmOBRwX5FQ7eh4aqkczet5xCiH0L
8twVtnCR1Gb8OwWfWTPOko7FvMNYXkv4fPkyrz+tSjHjh+3UGJ9L8tgLLHC4w1+493glicuCMXZt
+DHf+UGW11tWi7my8OhBdZjbmDzDkEs5huXPLKmKuNQL42a5D/9MOn1c7KJr4+3U3cFZPFcVo+UD
GRXBUxeTj2TnHzwzUMhFmpEiJGduQ2sNMOyLTUm0V2bPzTrwD9dsm26NYn3AD3VpH/0qkbPL2Jlm
Hzci3F6cHDFdecIFrxd8ZBFH2OWhPR/RJLuDVLQAL9YYtu85QCB8L28VZvfXii1FU1cq5Hdxb8Ci
jlHzN7hkoIyFGL5CSJa7r8i/efAtPwwjXUtNJR7cFUiqxY8oXMGnZQHF6GkBleCtF5dW18Yq9T3u
m23EWD2Y65nFQZRmkONzc1SJzDvqTrhgEhHJZhErDrVxpSYwDE1jWkP4mfoZnsoj2FzHWYcW7tzH
6zBZRqLwfoL22vrDbQ0jpbP6qUZY+1qG4YzdZQVuZx/ZswnfQpVvBOo2tnkNowB9vQnED/vERnYd
vKn+jHi1Kl0A+YDKJVQqp0+M0Pe1vLM0OjtDxi4quLngOnr5uzEKqdIicBaj62/79ily55uzd6gZ
G7Wz7HLCNYKNmG8q0+7tiWvIY3mBSD+1nGwDZ1wI6D0GOpQcCS6qzdi4aPc5zSTMf0nfe+KQVSSz
mg8IH6iHyQ54lfge8FE3f7flcblbrsJPWnQQ81Es7Q0HY4tbGYYd+GvnP37+i2HPtlmi9/VnbrY9
a6G2PlJTvn7lF//Z6aBuiQFUS7zBZleb06EYEprVHuk8GHD0alMTdj44YjUBp/0891s3kz3cH7ox
nvFlkevvF31PIlD5T43G1IPNqUJZbuEwHuu+fTAfMZG5oYP9oW6lTfoypKptk+u2gcqAXt8KzYc8
oZRdo/Mbr3FbD3ywYImX8x5QVEqHmyneOLGLLx5LmVd6PllXVi6E5gkzu/RQGJhdaItre+1eLv+M
p6dgp4gn3wxcOW4OxkvMjXDFZgFT/pCwB79c1VoSeFePlr2/4UX2sS7gMTyfv1SX2XEmJvvKVccE
ODwUUg2+Uo6tGOlFmvQLjOnhXDz1ct9ns0t4rfcf7Vh1N8hma7fSpw/NzmdMXE1bgUAYDqhFSatG
Dlo0aIj7iicQpklKFY3yUcA38FURtE2s5WGf5MJ4wW4C8jTYIKSOoNZmce9OcJfggRQSr+qSaS7C
bEGmwPUSEcObmLKR+AyofZBIdv81wcgZmV0rT9TRZus2rm4h93dR5WvWjKucbqBSW0mxMQuSNKnn
Z1PEfOUVKxK9cQzm+Aad7/dKvC5aoRIAzEEDqu9UJt6Ol3vu9gvGAuR79tkhGOINSnWUXkgQa1Hs
bI4/FGMwFM8pwk89VeKJOTGI2s8SJj4IxYyIc71xG8uyYM0g6AiCkFEMI7e3UiayTWxLuamlg/Sp
bNeQPS+e+OWDeztJ0oWM8SBnrLC6u1CU+XPu2cPPNU7c5SpV9IAEgbDKAAMhqde2Nb08/e0N5Spf
lHriNCTw/wz4Q3HtGdoYMoAL8gS+8O2BOjxvqAN8r+0g3Dorkw6KROBthtq3Np1XSuv/OLIevnyD
wDMjWWafj2YfEyJbZ0113BRhXJ6rGLI/CtgmIqq1nmzn+84g0A77ZZ0CHa24txpM89htTRPMnu4M
DD6D3ynI9QJzt13r/Q83ZZqWQrqFZb9uuePbjLI+Ls3CZf0O/oIvDMaYt2Z8z3jCYk5GVKPtLpJj
8QsaYzuymVq0ONcyud+J71BAu+lUbGaR2qQzbgjKsScyzF+gRdM9I1o6zeEmV5OnSG4VHXuGlHAA
wqtrJQe9TWKdrZ5hrJMRKHoW0nRvmiAPCT1JvlpcxfJWmrFY/jcnKMylYmhxkrCxLd1fRAPeATiz
EGuW5rvMv1ekatNAamFYi0+jQli1ogG+A0MXIWBX/hsup29NZf6T13fo+8my6pryHAA/c16kymQz
YquAaoKRvchEmsoR/18GWtOzWYUndFiRH4yIVQulLGUGOdiPxjyN5w9Gnuv2fLJQ+4yI+gMPxgkJ
cn7bWJrPmUrIzWKOw4bc8e5FCxPlxj4NnGcMr2kka0jxBcxiSl0YiUi3tgn8946Wm5OQwRmHmHo6
5sgCv790dEhv1E+s/HPFZkNAlnfx3o6wsuQ5lkru5cl7KUBzYtZMKa1ZsdXokU+fZl4+qJVO3QJp
XVjZvg6n1YC4i8Ng1OLKuwo6BSn0/SLk9uY6SMR+xL8pwwIycXsmnyUwAcnBZlhrZwWhuj5r50vZ
DdH8/wK8rTU7i/sYy+dz6bZ4WU0Ys4Umao7UWUODCoWFsQ8n3KvZMlq3PwAwkzO3l/GlVZWJs2+a
G7aT8MI3DhgFwd02qLRZt8uepM1+URskr/KUP0LtndyQsX8fY/ec9tJct3n8XIXxb9i8Wm1atAhv
OC/Ouh6BTSv2BYE+XeKYLYVwft+f2nzgz9ig3K9C3dBfhFb9Q3wHAhIs9zO0wgNYhLVmNxLaGzS7
q5PKrz2VQ7cJO3gflyWdxYuJPgdayXZ6/RSYvgaCE+N09KOKOECIr8qj/MIffb6jXZKjw1T5iEdz
ts7tZ6sGnpUmCb3mgKu6a/WgQq7HT1RD37heD3A3GNUHjtWZAmq0WUkAt00BTcuCowBeIa5KWrnw
ZUgGOg/ia1WCtPAH2U2qjEqliLW/BYRmQLNPWI7zap5QcLcDdJtOF2oXFGqgqKljAnfKFeEHknbA
huKxeIHHyc6jPAMYPNoZXv4DkNiV8HN5sMe7gXWmmIqkwbS+LiiiszB4rN1uTVSw8J7nblIG4y3C
BWUHe0JpxqOjha7ZmEN74GMkgoxazlFYqqTTKrY4DfyckKM0I4tOiBusKmF0Yl/lGaXS9f6pfptF
A0L4ghGw9tnCB1EG2yRNV+hF3R8oVrtKd8aW0LxgT+QaTnjMM523grK56Wu/xfJpoIp5rNN1KUd8
SKaK1lueuBMxcdcmMwo1Tewj6N3sI1tR6KVQskkB+BDpskn7Jwx0X1CaCznYTx6T7hH2arkJqsex
d+i60NHzVpW5RSHSj63c0C7BBodgejPR06AS2llg64YexmNU9B8hJ3DdMUc/f/qKm7kzMlVOV8sE
S770qeob0fUR7EYP/EU8q0Sd8FvBPaKrWYUIaHc4+ksBSWQP0wXruEbgAzLVwz0ofUFNs/q0TDZX
bOnUHYowbxR7xNF+kWbkjUyVfT3Ifk/aFYRVuOf3iQOs1NqHXvP9R9Tw2LgS//SK/LYWqccue+NR
RwKk1Nf7tPDOcG/rmIqZylDL5vmY79jwkxwlXXMOhIMgTA7NdM2MN8uHrKO0FBlvqINOqkoARyZe
/dBwbpNpqlNHriPvhXODb8QQYF5iKvK/4FAv9k3w356W74bpgWrqmGbre3Vx5Al9Tw9xmh8sfWh3
zVwGXB4Fdrl6UcvWaaXMoHc5Pu2yisycV06ZxQoKJJjsG94ge78mXx2ekuH6xb3TdibSuDF7mKyd
QxI6bl028+/tT1lAbdo/m1mjbhTkGTnLkq4KhmbCj2HlcF9BqbtR8H/9Da4AaZ+TKlpryp9Vjw+S
hB9W+YFUxEanfTKWFlKB6m8GQfA0yJ8W6zMs3c4V9zKUBxcmrqHJg3BrARUh9HeYwl+V0YB6nlPl
ORdL8zTGU4N+BEJJRquSZibCC1UaecYxg/ip8EJvoOBeKKW7+lyVKonB0NCJuzcSNy/JPuVomikC
XUbAGC2P51jaNTlapuBon4Uab2AZLo1giUw/DL66OqlGaRwWZWzgrIBwonDe7liGQgZIdBTQ1/+m
tkVBdgks2CYZUgJvN1UAOmb4fQ2StOEJIxiwgGKgeuWfhFmOePhG3Nnh/AxZCXK6gkBcvyUQaQDK
UGnbrY1DJ00OlISe9R0DKWDIsLSHaWfwc3GS3tdPxoJawcHXvLup/S4EgVCk5LS6GMLI+t6cMrEc
sozaq78YbTT9v10uKVuOxRQBITLYqq3qaPE8lif32rQH3NQOgaSVL+fSsSWu4BVZuNbuAu6IfVl4
cIJfV7p6i+BmzurNhddV+tdjcSpCXODC4wyVvLNoH146qnMjFMkyeb40bOjQ5N1PMzDupkoc/hLN
DxshOWzUGSEJNQULLspq62il0GMERXKpqszT5F3JneUaAoT5sBQgv2vpGFP7zcJk/5qq7Wiuox3w
3eXXPbcojfKKJC3uQQFyLkGpGdSIt6iv4orC2QBjU7MdA4XTdJ3mzfOvvK0Q2LO5/hmwksmsB74j
wrqIWxadyalECoALlQmLy8x0JATbTiKH8J9m8Ik7WGg8zVIabmPDy7wxHqTIsrmQt/TTDg+FOCNd
jqgIS9P9JNXKt2ZExPX7QGSYrmnoignLFA2RQsf/ZC+9Qvd/ZCNtmNRNOKHDJtQGzGJU0ebLl0j3
pU2FCiM8MKiGYoa20dthNMcI/PhlGGEK1r3BZeIYHPaHeOt1+/6Rd8U5cgzgVQ0gVfIa48Mty3/g
zbsciXI/fhaTAxvSRw18Xcfd1i+YLzNZlniD1atbpHRxs8m3ftr750NMsQlcgBZrQkQe6/N8EtYF
O5dAFaIHaWX/UGWq/Fic2vQOdVJfNkO0r9fjHusBDnNhtFaqrxzvmmW7H2bK7JGVYzy6fwCEex5b
wolqvoN/bn88rXsfaAykRN12V4l439def2YDO+PJvqrWs4iAsoavUrykDiaT+vNkU2xVvmQUpCqC
n7JnkZdRHgMeSH0dCMxvONuOI42nXmILbpzi9FEpyZt6fGYEgq5/aTfZMC1h5BlBqXiwKs0Q6GjN
bmha0c+4Qg2dd2uvDWdRIt6ZDhiXnJAMksnL5tAqYny58xBzF8SgEy03MpLX7WRLBN/axUCVWohl
yugd52p5xmmoEaukR3dBTXoM413r4PbH3Q9THrrlo0f2Xm4OMSCmJD8TX1GGO9OO7VES/4H5WrPK
qMbauLrdi3v06sqhkyRlob44dNx5RPX32+4dKQIrU6hErhYmOiqeAwoGipugCqUHqkuJI/NxcMUb
0sTmuBkSZBf/WMCfv66B0lnuEIXdtwWLsf/dLInFzmVofJU1H/a346icwlCWxXP2M9X7tvIO7a9h
8WrRrJjoqt07n+msxOWvkmCGs7OKoO46WZO2TG/95SRvj/eHwPgTaUI1tzS4t5snIcljVvuJEcGe
+6ZgBPN0ra2BP1GnMk/s9zhKeSvpO1MDWDGZvxudQ/msjcSH0P7uxcU/KckjnLKa7AJXwmbP+WVQ
cOTKunmteeUXw83FoBqcuxt2DPEdLkcIWmLBlDvUalZQ3cArkvkIBVoW6yEm0TaTMAEdmi+FhpkU
LvH+7cjMEgS7DsbyVARpJBJluG0H9UESss2Ccjr1zuElI+CDy6/YqS8pmxL/yySy/aTAZbqISuB/
GV6r/If18quD26pI43Un2yildV0B3MOI9RFokx8FbkrG47DeWGPCS4FFUgbuGEk7+/4kzFMWw3UK
4qFgn2VvyXfPwueCaBeYcY5HxrHVwL2GgV7YKf3TjvSrcXv5Df9t4LKiJcL6u59dNw8fLOv/ktSi
Vng4mOM28nM7aIluaCJzBbK9bt1qqSB7eyDlNPIKugRCMO/gn+p8FN9fRx2Iyhi6QA8OH3KhUiG8
izAFiV/qVUg0tdbz0b+Yftq0vdJUycLdiEU3mWx4JGnTO6rgCynNQQyCbYN3HjoqPGwgUvAHtbaz
eoyNGNItlmkOY8cs8bw8v3sG5rGlDJrGY28fgy4xZZTARmXFJpQPVA6h/M35QQ4h3yNBhXc+bwu8
oVQ8l76yhzLEqzsXfApV/DldUZ5bO7dtyHn56jPUYr+9Ze5IE8ixFUqFkKThcH8JqCXBsZloOtb9
nFaYfdNB2VHZFOMqoAexj3MCUlIQuEVSsm85orGJytMiHykknoFSed5HZnF9E/idWv5HT4RJ+ILv
6CGJwGEU7EGzZEH3pJSH7mh0JSW/Vs5OaroQtI2MMR8nLl1r357k8MZcz0TPoKvzp84EXF1eH2mV
Liezn9RVqCrTuAGwMm851roj/oBIB2nkAuAVKGoQYXSwwQ3SdHTCvLGE/5aacNvQ81b7Roddxo8A
f/RlMB9YD0TFuvZZjfEOhWAnr6/oNjdq9/XOK334cbPujSMKLIm177sHKfVZnzSEGHaiZqrOwiuu
YzwkxNVXYDqk8ufiRYm8Ef1horl9gAI6UgQI09MyYup5B5SRixMstOxCd+w9a4TPYC/vSj05U5qk
1nM7x82wpd3BPx3PmYf6on3R1lfcqPTEkGDx683KLsBaMV8vDll9hsqUDbEUqcd+kZXsjJky33b6
9kkGy1kxXtYBQLqor4WQ/PpKJEuTul/hwZESbPcIYwxLiarVG4SZQN6o3oincgUU5d90OCPFkJXn
XO9n6JdfMFiVhBVaCAwtNyfGin6jaizBiRRZmlG0misEzbjMTcbhEr2CAQGoyKTyaveUMHkrjpiy
D33MT4AwGQRnsNhcxun5Iz5Y3V5+Bj7TMlbc3DB2p1PR6/sNhn3fi+2iVznkOm3wbKig+mO9Mjd8
BKDl27tfY3811C+FBVshGvB5TMY15CM9flt7OM0LDMtb0HkfxtkOmrqXmAM3vQDX1OucpqD6Y+s1
N9oK2f4qyJYONTTy+qPKpBp0SEnOHSBTgjhenZwoEWJMjsB+l0pFNTQzYOesTYSyOxyE9ZiJgRLt
TVvoSwCeMMizn3PFUsrgmEeF6cZOoaznfmNvgPtQlPSY5pUzyFeT7fK+m+GeQx3ZM4O8iyHYMiQo
vMs7fEeZ6NkoVf9oCAen9uNtRaym3RgW7gEIDg+XtqxlmGHGfbb230jm7z3WhoSiWdGxMpo1c1US
JhlNXA6dbnx1C4F2tBp12MI3OQqvdUuXeORhZqKJuFLkgjJ0ImAeqjZ3rz3NAafaMY5ZxwLqZhzq
cNuwaEXuhlu8/TP5Uce/Sy4KxG2tjaWWz+w/sSykjawsQZXAeV6WrLU0L8psUI9BH4+6neqsWe/x
03jvP79dKqAEPcoXfb4HsT8qOcUWlXuO3BvB5Y1d9HMffMcluEA7ojRsxE849kwysg1YC6eMksGP
U4ssu44kcsbhDLK6dm78w6C0yHd6RKAoqOdkDmdZFt72TL2RfKnCVDudrcdISeoPFw7U5odfUa6+
b0RqfgzB9eOQ7McRZcjEVJxdvJ2CKocJohh3IfRWI2GUXSDYH/+EWw8l65vuKLH0Kkb8h42hLNso
nDlIpI5JYfHkxQJmAPrBC4GQxlY1rNiG2GeJxZ63hBHPvp0mUJcrQDqbpUzgEX00EYDa5NSFru0w
Kl3aMSDRjxzpOjoe3uORp10bPOuWvk+jP6j+nFKG5eoECgU63Wk1mEJKs+10RynPKZtw6u7XFhfP
jAf0yc1GOSQfq6p1Zsv10RQH1qChiPy8k1iyyylLk9FhsIkrVqZylE7CHG4tqL7OCDHN5kGF2Tg8
BluuqPt5BtfykCs1tXjh4CFu8FYqfnup7c5BSZ1hKyjaNqoHDHsOzIVd+eFGkGLx0osQmSINC3S4
ROdvKb3H1bNuR05C00ew9Uny1EYlhIUMDCFlbzh6oBQII2KTQsd8YXudzAdHYi0rZvE2MM5otiAz
Roe1o2OzuyntrUoPBQA6IyJ51Z7EnGm31LTJfSNvUr3cr6300ha8M9H56MR4LsEg7XgQ6u2uTD3s
RY0FDGuVhR6f0CwB8SnY95++ejc+UTT5m+XkVCqNbZ/psispt7Gxch4wJ0/GvrXr+2H+9kS25BHt
5pNAYOrcyNjjo+US/CTqkJ9v3gvjHUzt1hdkv3skRC8dG9fgWKwFjV45mDHWKxHYPsQLHxnsVqfw
vPiD5QXEwwyQ+pz0h4nU+6+XB7qFqzYqoscu3WvAGov+VL8z6y2lQu2CKOaGxzXdG5v/TSnt17Io
+cqKkxLdLdUEoz+RtRWt86qrJbXQTZL8QGKBjWZ5Jmz9T+PngxgBxhG1CqUZQ5IWKdwCn5GggmBS
FnAgW4U35F8GiCcYDsVsC5kAAQAbg+8M/cGKE5t+aIw9+6C2zyDHvrGOzFTMtjccS1ge+WHEs+7T
jZup+xPd7r2Bxhn608n8PlKrWTItCA8H2FcbrVt891ybq/FjJMEEwvRQvKclXp0RT10lHRzqQKJk
kG6xj+n/vKYxx0gXNkQwGFhFRwKCiglC5cqiVYFhGLoj40hT9A2mmOs0/bsP7I4319MwcjddTMAW
vPC2LLGfsvJYLhnKkTjczMb3i9UiluPMC1zfTCaGNZpxlwxcpKhXYEMuBPgaRqtndQVbw3Gl+6Mx
ArrD7Eb2DCYzFUG0tmQbgZT8mrVQvCWGzLMelk+WZvcJeS2l5mVS7ezBQR33H72UtaGUoB01jb6J
n0CF5lOasZo10+CPPpQk4CR0k2FINX0K+4D3oC1Hta6Lg+L4r15ppZiL85ifyq04sp1ttVKXnZoj
24Nrfc7NfA6GWkr7quCwBtDPkZiYAt19vW6oSgxbH9BLfeXEpQJwyCsN6ozO5Lz68crKD2CADD21
ErjMaq6qUkgRCpgPK1ESfX9QJindea6rXwMT8tQOrmb8UB0W3XgBKIykWNOzL1mdfbKgXzRw3osM
rYVVO5pDMQWC778FEELLPtiGu4rGGtAG2/gInGQG2BEZmNbGmyBloLKR7pAzWIk1iGhR4Gb3q+iz
nyIi9o+l9hgt6p0Tzhh3UZFInsigSrmtVKjl6g5aUbkUVwDwfxi16Qf1pBb9a23/oGulIedATRVu
GipFi1ceu8WjLG2HFCnk9b9C4Y0/SK7bVw4VJurfUYhRDuCi70wptw8FfptO+ik3NqPPOBYcHaSC
GP05mo70aDcHa3isnzan2jlg5ovo9JZTwjLvRa94AwZKaeqFQlndkUet+f/tRcYcp825/kcYHhG3
FJlDKBecWDLPPI1RhpOi49gRMYHnX3Tio9U+LgIEEtjSIOm2FVmzQ7vsH/R+H2ey7JhpC8KQG55P
Xel68BJ8G913RbGwMIUSCOuQAX9WsWNayiN9s+hkMxe8CXwyywjCXoLHweSoy9rOtqeclWgn/d1d
6Dp8gTHsTBYEclNWuX2dx6j9CxUIl5RBjRMana2ZxhnjRpmBSCvYceL3SYM2LUOXv8DAozOFH3e/
L7mEKTAC6c4DjgRlM1HSyJPHhsvu852FFpSJM1JE3JqCz/AKIeKS5b9hDJVbrhFWKuoUljFdhmVz
qp1NFHRuZ8G6aP/MKPnxYsgPoN6TYyOduwBQHHXMANv8ce0HlpzKHAorrRW+GJajZlElS9fa4Emq
SJjixUNSkXxlfChsycgcC5F//rVtD5Lb0GZvOihk7BTK2mdgDU95w2XcDXpeN6bK0f/1wxXtVF3b
5y+vEg2pM6FMUUMVRN8xUs6a4ZUwKB3i0O1fesM7zIAvNNV7gNAJYQ5+yMWb4oqkVxSfn113qBMY
EG1FrOuy1o5Vh4Rm+xUh2AUWilmcVBwhcifqPHcLMRFn0Kh2TK2v2EA5NOdXamhvc0H/pStZxtzl
VJijp4I5w3uF3dzAAQcowINKXHhoSgAAlOPxkcFzH4EoHaky6MbRNoOD2Q112o4/+WVvJR2qf/Ai
nxZ6d2lyFonaC/SwKWHwH+bbnb6aoDZbxNs9g0fMzJevoF9ewgOx4UVa1ySkaqaTRidb8kWljmVw
/IUxeqYxrWSqXm4MZD28QC0QqtliTOlz1qPCz7dTDhbr3J9H7qiFzcJhhTUkRXm+1EmN5ar5xlrr
jundwY6jrgMqxEAXMq48c/qgGRu1APE1Nr8eReTtPcTntwzyc0gftDl03O/DOX+XiFN9CzfALaCv
W1VBWmcc/9baov5+Kq5GE5RetLGQ23597P0Yt8oRu3DlWnyXmKyHOAYGqW87c2fTZp7WOGD01183
ANgM0d131aj7v7Nqgtq96Yq2xjKEJ2r8wJTeQiEHT+xR+5/GTpj0i06Fu2W17LtCSkfrflPQXG9e
JedTjHBEANmfZ1lqRHV6M6eWnZbmYl0maFTMfyPj3hIyQmBAONuT2A8ZG6eNxn9lDaL8ed7IwlDO
iWBfu/pyHgZcnb/KgCFH7NCzgec2kIq2WC/y/kiH/8wlalyySZ3YgvWxeGRCEEO0ZJ2b0eYdkPW1
NXLPNUGrbMx1ywwWwAcADKRmYk8nSFV0feL2JiY7Rz5OYx9lV6uKGwWq8nis1M2dHoc1ZE+8DQJK
ucO58hjlgTMs02h/rSUIGTXtUfdmsuDuanAdXzH6Aj7AEzxBq4NXkTF9nJ9+vZB0i7hjoF8KY0AC
yR0wyj3xLUs5GaQrEN7YIixHHg5kDgoSayttsdp0L+vsJpuaBXSpWv0sUAYdOQOHmUwsobLn9ED7
7H4BSuSwA4eFCUqe/hApCyeXJEhuj2v+HhNEcHDFh9M85+dx2eZ1PAExx+VDhIcFwFGO3nI06bJ/
4MykpTGJE7cHTBPtHnugw8GP9khKVnxn90VxXzNWTFcTo0iXe1SfM9TBqMPbKoAfNRx38n8MdOFm
S/6HbFx4XgAxyD2A0m4gq42C53feratoLUyTLGYcex+U/B86cAHzN/7kNElbkq3MnkluVF+B2GN+
e9oz1Sl7nR8S/Ythbqb5ggcMCV+63HrZjxPxMmPcbPJkGoj66xD8cFvTs/iHbP9xjIaEeUeyGVK1
1P+GR2F6sVmaLAKi9tJXYyOh5FICKkTQTp9vxjdw/aNhbHzYDJ6T0uIWDGwxV+WhkmdWVJfjB7Gz
rp/u2bnu90LzEx1WR0bU/whwI5ikFT2jBj9GUXeBez0S4JpzMfIOfYoI792NzaoamAvYPGqJahu6
mzx7zaQBOLdCadVkwiVzeanhhyKQDR7QMZgbg6HXa1AGfgMWp1KvH9fOclHskzLP9iiXEBiq9dr8
sjmbuD0XSv2o7dJjmMlXcj60lICZo8rdqBNoDG2yj/9OW9ZTl1+baXqI7M6ctIpetv5HXeSorxeF
bd+UoJoaNjaWsvmVNXLhkUIfCy14GxBaz0w7GEhkSiTg+nyR4iKCLtLmnrRnmXLh75dRMuk/mMWi
+b8vP4w/PN0RQQdf9KQhQSxDs2yg/FXF0wIhR1QkU+tI8DtXaoXD1Pziiudw2rdM5jtSglnfsI8f
gttRfUQx4HnsqVWEJh7y7Uc4gFCt1FS1eLFzK3QJp2H0uo767f/un7H8T2YHTWajCP6sSktxakc5
fefWo1RJoemEa0FjglfQ/iSPhgofjZjz9pUEueIbIiNsnq9omOcqeCVXHt9C7evr++c+UJQQVnN2
ggx8TPPgHeSTrqEOnHpodUgUuGIUaWLmVlyMLWMm+A+gdVt8+u/1nA0xaz+d0cqsZbapVn0W/w58
MJIQfNjMDtcWuRZ2vGNsQ/Cj2PaJyhiBsZ4umQlssTl+GxM66YCLRIqpe8v5yrD57LesIuInfNlU
ONlnAF4tHMPVoeiG0PxLVRbCO4Z0COb3MHUI40k5BTVhvCgMsqdZn6rOgYg57tcI8oBWZX37KuT4
0LYBAGKcEkN6eSVEIMfK16NNpLLa9B31wKOftoUf1RMmmcwoWRk6zTzB2dkCi552K+ULy629xDui
iy58wD2axWdXtVWn5d236/IXJ8YV7lLSLC8g/RZCMZHYeH6Xk4CaZFrtjLE4ANcZMK4sTBPCvkTn
RzAkxu4ipdnLabrgBm0ELpQT7qDCiTUsjLWqSpSULFWHz0eT2ESsh30DFqqFdFup3o2eQmVTZ+Ka
iHsIowJkJWJvqoOrLgjK/uD7Bf8s4WPjyvdwBypfS92EY2iAyqDvADD7xTNs7eCzRzlibHYe9a83
ujx2LYdcesgypyawkscqlw9Y8r1TyF6XouAY0MXfz9urf+0Eryj3Buk+9YJ9Xopc26wUmmRA7KV5
MtkD9gDjzw9E29rZMbR3mVDBIie/CpwFWYfmG6sgOEfQmvdapRyqvbC5jT5zzq7do8wHLXaF1GbU
mhzGczGm8RsKAzpLz5ho1M7hJr+y8CnUTsdwFNUghtysk6xkclT91yuoz8MuBDueIbOU8E1oXFxw
VS8elT7WCvvYYBiOJX0LQGrQBPgk2TM1fR39W6zFA9WR7GioziytWNJ+TE0CED8lzxmpbtjeauhu
9038UmWyTguVq/kYcsC2zENBwdN9OWbfbZFSyMLm9q6hLXdv/mVLWppTlUCm3uq4FNYVFEhA50Ro
hiObyDvuSUDx8tM5JYpR4Y9bSxCUXKIu1xBJ5EunI1ZhYapMGB+MX+FLzOEPOHOqYPAtTD3CrDR4
PA7ZIz1C9Unj7pPTpfA+PJ62QPldlenBF3r4J7bQejrsPHekoP12Nq0rL08odQLDpLi3cHgWRqDB
1UfnceuCG1Fqqi/3UM6MLz6/nLn+VrwCNPK/H42UKu43kmGrp15LU8wScvXuPqbGf/42C2RTTJ+t
jqzBkykJ0+MPyfBhVo1pPQueoQ/bPUaelwafCDhUYl8vqdvj7jwN9RI2I9HH41rzR2LPD2O1N46j
8OL6Oumoj2ZWd+bPLMD3cNRvhjd2JY/XpPiVIp+bisHTEQi6vk29U4s+iKrMy6/2uPS2UlSwjPOo
Hja1tRcFzyJBTjxQf8rkamH7l/ICXFzhQ5UgaSXhjQb1IejCTpmVbpjq/xRfADzgpvJSaKgw8xPt
lM8vf6kQJhKwxTXE4IV+emPugJvRFymvF7YdEQLWypithct1AXs/O6NwrXD/iHwUTyIKQOdxS+fk
M19kSUYH2aw5PbXl4MzqXnPdozF/4EuPhYpoFrCboBnB2aM9ViMi7e5PfEb2foecDM+Kr5EftcwM
7cYoX7zDoqEuRRneNez5C9NysN7eoHjmKLC5QXgSp42QzR8znYwThkVGFh9aYz7IbowOOjkw5Ehj
LXAbjPTqs5Dgpv9KYm/OYb6c6V0sz74isG+I72ukKHAfjXANeMcK8Dqdew5kk1MsSRdkoQM1pcWX
wT0nwO5KXo+to7eTtzKhU0yHsYf7JnySsP1guk8kyyA5RWs0CM0w0i260/OoQlMq6gAvCtnxevgO
HnL6hx0bkXN8KhePW/a9NHqvCwvFng84WO+FW5djGvVVjFgczKMLzEFvSqQoN64zQ8ZXXxKO/CE7
LKsW07uIGjCn4EO69v9SIbgBNSmf6+TQWLX0se8yEh3rzCP/63OST+/RJS+N+xJ5qUUZABBiIxMS
DnkGHdYH1788iw9lR3Z4Pni/hTm1Vy9Mdl2J0K784DZ4laadHX8N8GYTHlVc7c98s0k5ViG+VIba
i4yaQjEoseif6683hgMWTRw0HST2t5Q2ILhKDxtxr8cY75yEHS0kGKc/7sxtfnCPch9oD3Lktg5R
wZXcaJoHOEVCux+5xlIA2WGv+myH/81s5GDoV8zA0IRlWygXtO5Jol1CbZGp3YauZResdWY01zuS
4sJuO71dbjRzodevHdw2jXv1OTRcWHZmE5/uyJaERjhc3KLLK3aEOXCCiCYV1Mmr2Uy/qIDl/IMw
E7Fj7DEIWIry5XvH6RmXvzUoHPUc8RawX+1A7OWU8DJ9uNJm6EvpUWJwElBeQr+x8SDj/1+E5BB8
LIpRLMlRWoVRvk3bY90YJjYb4G52Du+1+mSHpgd7ruMQyG5MHzIfbbOSukEjxtYOGOzaPYJwIKSP
u7C6Ixw7pBDzteawe3c1HduNCNAxaqCr+EkktP9mwj6WxuosHfuq2JiryIFOWWHrcZz6LhXdaAmb
/G7ufz7i2XiGZriWcCMToIlH6MStGcM2DhKM/o5Dfi6Lr0U3JBnEV/Xr159E11P6C3eiwIL0KErg
lLXPplbvnhcUPmTebdHta9b4xIdQiQutk5SZ/okCNfNmyc/Y0Z7vRSkEomXvVkJ4cDcP61ClFhu/
KUWfv536CpeM+2xmbQUJIQ7ka9WJGFnZGppatWfy49LmZBBxJJJQOjL7waH7BCulmfxMYshmJh7l
TKVgxs/37uOhQbOm0Eo6SfR3BYi2bCY9Bdt2nrD9CC45IwKjf/ZhcG79pxSt4yPVeNI3PhvJKEdI
grKnliE4M02HHfbJfByKy3cS8AGw6j2wLCeNV6KBZPJkqfW5dHV8fbFjyCuU7oz7/RD6SYir+UMD
c1CAsbb6Rd+hbo1Nzx7ZZDUeLzYbYf0jqRzCYR0xvk/RcVM3UUQMUJqqs2CKVLwmg0fdbgeN0FGL
cKBZKUb36eYwc6pTil32PVce+Pezm6DuNhjYIN4GOFcsRtSO6UZ96UqlVcSL542/sTpazxnNhm1F
v8b6zsaCcGMMLL4xgzPcOeq2nMBgwnsA4IlqY5uOSET+621WcY1ma3I88S40IrwY8VCqugzRBywc
f1GZD4LsP29wWtjHJh9soaG+4NRj9zjCrLhLlZLv9wH3G5ic16pEvqTvIMuCEWRShsGviFG5qqjk
hP5rxCPuMXjmlQtrWkgrmafFsGJqDSYMitS00WLqOGEHOjIkCBWAm8meLGINg6QdlT7zoozaEjFb
d8mdLBtte0FeiJDXm07dGW+6WRpPtx03UazoCjs01L/iIpWfIT+NoAoHpO2cQWgsGpZi0TcND3IY
AoyZepCiYeBnlBomRPcqcEgL26RXg1I88J1aY1R0L31L2skxbcCN+gQh3HWznpF0qVnC8C692Mpy
xmsEen7dy3tk8KXpzmNtty8EUhexg6PgWPX/TRkCPhmAvbzCT9XyQuCQk7x40gqqeT2xS059vzbS
CLn2RFhRR1Uqage0yr3XtPpgFME1wBN7kvMqdO7HY9SL6DDULVWGdoCNivpsbv3Jl891yxzJl+pq
ozRmGp7JxJkgfhs8eTY0BYI+SnRh2z/ey9n9Ccy76sbSDRFpoGqdtn2h63MugY9yHwqIn8V6fq0g
kNM3ncTwRMCGwZysdvp1KzBPudIHonT4uU5spnun2KIalC3ennWuuuWVEnvdW216ZRkZ4mop02tD
GMOQ4a2mH3emrXeICyEtho8oG2dtWDA75Fc3YnBwZoqLAHwKYvX0UtNKdnEeTNayYPa4WX4biR1R
eLxyOi0xMysiFXe0ik0i1w5jBOIw/DVPeE8Sgohre9xB0MwsCJsLMFotcLNx5PBTzc/i1QBgcAwu
rquvILG/FGfdW6kmEDKiqq8ZOLk1ob8Pk4UpSgW6MeNabB538cstuX/CH/LAbUfClhQImQ7fnTD0
pLCdLRbUYISmGwUM2T/MDPBmvZ4Ve+1t+agWKbK7luE6BW138/cWG0jRHv+aMBHrbQKgPtQon/Uh
gIjP9erJCv4eKQgntzNx9xm2oXVaJQ8Y0yAhBSKwKYpzMB5m2pRc2cABT8VJQd8Bvk4Y+BjBAw11
wWiTu/Wq0HfzqIT6edvxOD4JnxhCPIGRIiMWKx+kmdegpyzdVpN23lcVR32/T0fYf/IgjeDiS6PI
qz2hPdALisPgzCzMmKMFrN8Dv/TRcj8Ab8ZZKBYsBLuHqdMT9dY/pKtxZ9jtQ6kzaNCpflTJ0Rug
T4iCgeYkP7/Umvto0igU/RbDnAWFEAypLWEgZA+nzHlNBJbC5BxRJ1tZXRTI/bua36EHNQIXPHs9
xbo+lgLFI7GucydB1gfn4RGZckE2vUfDcdyEIM7VwF0c66n9+L8ZZvC8gqFhTC0c///lMFQP080F
tMdBvq9YAimBCrXyqN1SH7s8qL2Jptlc1xhjgUaw0LrQuDHKVmcq1D0cEWqL4b3QLf7/Cc7+7koD
QXceIgBuqKqanP6SDq7H5P7TEaL39cOLp51KwpOgkeI8zpLZc0ma86O+dkF678nRnKmAvhp/Yub/
n75ADpo/VJngW3FWJt6CodtNrKxTF4/ScE3bscM1gbvIQUSBj+DtyX4mOWQSvm1Z2RKbvQaCzqvw
JXsDE1ZejzXiVJN2y5C5lc1Mp9XtHOsnQ2jDFFN3nHlRy8WFaDWBC4FzPs2n0wwL1oROw8zNywg9
eRDgrWb4nKr9MKNWRb3sIvzsQeQ7Hp5ST/mZ8J2ULqkMCjcYORD5lM5MX1C63yoavYbRccFAqkHb
LJAgBxMMteVjVCAZNC4W6h+GXeitp8uG65cSiipxQyB0RRp5GJXw5+Hd/wBoaRaHLC6bq58N2KAh
Elkvwel2P2CujL77qLSlESR+yVbg6BVFS9elQkmMrtvHEAQONUpaL9s5UhiEMausQvBchRN6t6q3
oomx7mJnXugtab2FGR0gSzvS23vhlVfHaEOKa02rfB48yGsVQUiBVbnc4vfOgScm6y8/MpYZlNny
MncB9qP/KUDNT3qUO9RVRSDZnVhbDLN1RpmLKj4TkdxVqsaq98DB+gdSLN7SkBpkvaYL4jCpqHuG
N8kHc5DrpnnD724T8HXHFiIGqjFFe1wsF/KyY/RwOiEI60GJ+4Csewlk6PGoL6/Bt5SvbJB2PH+o
8Uh4hLIefBPEIrVX3xppQsUKcd/+aD5SyzxNEaXcLM6ObUQbhpd9RKiXgCFPHsbnphNpSGDUSmm/
2d2cmhTxTIdRYNOnh8niPhXMWkFsiOQbhzoVV25vmI0kYMAho69bO5hLNDKE4JMVYrUuv7tHLcuj
f9k+tgPjSgyroT/ZZHhq3kOSYT7jcmHzFGBUafOsltAhw6wxv5hwGrSQV261joAFpJS8s0UW36Ya
2UJusNLiVAV/gv8GgzqJPNFg25KwVU3cyR8IrW9qSwGx6vdx72L4ropNRJ7lw2fys/wS7kScKA1w
TQxouzstaiUFCLBvhduux7dqCWjMjcV0Y9d1feqKh9UIKLzUREAUxq1TmaKYMMBfxJM3N5dHTjxp
YC73xCxcKYlj2QBTK4hg8OGg0wHP212s4lnPmX7b/0AgSqZhkb8QIxFd0/wuOeF6z+eSShXs6W0Z
ctNMlWeTQXfkcE9kK2P/aG/zQ1yMnPhz3ANh0yIkPHBL1UEehe4gmh6jjgF+8Hh8YVam3fpOS7qQ
HxXnCWPVoo+Fz7pXKI9SaQuZMdU3cxeEmzEwDGq05WA1GW6kKJPAwRFPZINedSkmaf71GJo3T4bs
cfuAPlYKVUoDEg7ETZIeguaxSYuG2y6PcXwQgU9uOQikdKKKCOP8lAr1sNoaO/1u+2prZtlbUETf
NYbnxB7x+8dd/ewKor/LHcRXiXbYCgfYpPt+7q/vrsrkBmgho1OnuUWeRSwaq1a/ugs3tx5K6IR0
4FBtvNgByYIe5sFQ1Giuhyhyf36sECTHxO9raoZIc4e5KgXm1PiF6SOZUbZVEZa7iCddLTY/Zkfx
5TW9NQUDWwj7TTbX4XlxTKYxcWLF0JJgbCU6yNVYaRO3oxSfqw/YzI5ZJkd9xQyzSfVbVHLhTU+i
INzM4YRZyhhARA+o5r8o2zQV49WjsKVentkTlWTONpahHixyhLhWEKJkcpRdPbw4fE2tYj4ctexN
ijl3mGfbxIm8AVtS2BTg2Ik6JxtAa1J3dG97ON00932/JIIC66P6+vOOkImUq62Yn9GKhzD0Ym0H
KtCi9wChbrqbH+0xudT20vCYK2QX1nstaMAa5UcTE9Mr8R2ZfMQlfmxK2IF/1Vks0TIDTaO7pkM2
qo3DBvMm4JLdIPCXkD1ng+Aoxfi4hU7qyqZzeecKgx1EOy1ZQcTY9WFMZHGHKUTx88Obcv9Mx/76
hQx2Pxi9m8losym49VFA9mpWXAJSAtbwkZX91SAl4y3HKXUIwoHLL2C0Jj4LSv8yFyKvvi5rcRV2
E3VBBehkwnUhvRVJFpyAsraUKj/gvM3tiEc8bvOmaZhdcN4kM1iESKCXtoODaCzlf7O3mD+2a49I
sfkObSnIUzIubmno4XnHB7IDC+jHboKvlNOZYmji2zJJcUer43sgGYqzS11g3KgkAtCf1Y3Urj3I
IzQXlCbLZnOztje8bu0/TvXKopRXOgdC68YQ1X35v9JhdoKPX54l+kkSBDAgtalho6+Mzd5Q92DD
EuoLRU9b1Rbehd2eQ9dg0wtGh7TgEqbX/rrc0IErsJukt/G5e2hIZ+mTSJsG9V8VvpWSA1t+HxZJ
v0HoQ2jKoJ2I11C+g1bV9bIxL6Tcp3GNoOjzzKuSzD788jHuYu9QgWboVN0/dQVtIEbf8Sf0fDkz
z1/iS+wL6LB30gCD28MsKrIvtjc56X26wisfybhxq6qhCwfFqWohNUdE23Xygejf+c/yQLC38Y0u
K8wnJVEWHZUKpTsF9Cl6ZgyfNelV3zP3h8uv+wECB20bLdlA7lbjlMUB3BuTSFcNX36rgzLg5Mqk
pMY1849Rnak6fn67jiAnTb4FamBgkf+BootkPXO8ELCreuhoyeHTxjK0TSqxalb3+/N4t2PptFcs
wNoodiEHm85BYfpXUggq5kXKa5en9hTcHTppb4vXQ4hZk789obx5Mv0CprMiMr2slmthX4GYJysf
ipeRZjm+He2kErxL7T/jHicBnMvJJgo5lq7/sV7uOJIp59FKFZDE5ZuX6N6nosoVnNmO9DNYL8Lo
NnfbUlW6Wc5Xhkj6srHO4Te2FgM0bXJaFIMbPxYBw7F7ZpzC3INOqbq1ev8wvX16EiKH71NB1Sal
f5SC2AzMDu2WSAEF0xVVby4P03q73i9r6DJI4oStk/2nFvNsI/wc5xhLOobErE+hS8nLdJOoMe6Y
mBJNL8Zw8EBmhKhAiqmjcetVLyEPA0K5h44WSvKFgjpRXozxkHaZTIvxPbOydZaww1z/b103ReGQ
KxtdDVhUz/2tXhdHz/z3riYU8xwtb0cFeOe+2NeuLA1cUCdlwbDNmyOCmnQz0ii7Ga65fW34VKl9
VsZSw8difQ/x59Ri5v3YXYrJP9eoGFh954ZMOUgOGjo5SUERRumXIkVxELe0vIkYTrWOI+WLr/hd
4RqPPsJZ45uN3SHFHjQiclG5C/cg70vVXa9N9sjon3R7kaxYZq60ChSf04qjBTHr1sGbYPQ2Tepc
T2Xr7GQFhKLrcVg4nM1lfGdL3Q5hpkhMCddLW8KC08QYndOZKEssRWPtRIP30a5r8ASmeK+UxdZt
E8G5OEAvlydTWzhmGU+i3jc5ND8bowfNjuy3cq9pqHZvA4G8AbqSOE1WMZqmqa8wr2RpFm2xDS3w
O9Wi4WiL5Et2UbUdOD4B2WFYnjQVYXtkrRrbw2fo3KvJaTz7zQwhuKRHednl/ve1Mo16MLZ5xNdq
r7AO5vn8Cw28a+VXNoMEWUARX2N1KpFwsTBGcgfL2AUdgL8+5QKhG2ejX2SOsBgj3qOABG39XWvA
uQjY1B+MtEzUpiPvUe2O3ljMENaEEhxwzubrso/oV/gtDTK7VT+tt3MJqNb78/OMeuAhDX8QfB/G
OVepPS3RR4Rf+sGql7JixYSGQOlvpcSqRhxFwDEGsR+9nZgdDdKbM2PrTXOun8OBrzxBjqUPHbk8
Jz/KIdloXoCDm1WNVf2JI1lV9JZoG7gLIcHCLSCyxN0PoWK3lt0bdwEQ3ApdUoNxWbGPR4+nSVfo
HR7hbiCE4V//3C9Qb0sMenXCCmPkfsez/kmO5iy5fsiHBjaogecof8E7qbXG5icwNc35VlVFxopQ
m3zRuXB9FvYXPxxMFVAcTv2zx95STcXg7oDabgmi0wRh0X1f8PbwlxlVnjINTybTtPn3wL1m/4Xx
Y7JHevj641qDbQww+5Ydb6EzsAwsEEBH3HMv/lu+ZUbqrdnKnllnNcPwT64RVmiccdywgn4tZegz
F8l/AxOq6kguDJQOBk+ofKY6Wj5JS34VMdu40Z59odCRiNtzV0sUYeUItkVNXHPcamslOWYEGwrM
RbKzw6c/TywHU9W8dtt24DV/b+nSTNtsAzfUCohy316WtfMdK+jboQSET5D8szpW5Z6GLFQOn8K4
1FNtN38NXg3IXhoqlf2G3oDQHLzQ4CNqYs1M0oT4y6xEtgilUxWxkbQaOv4/4qRB7sgpPnzUgEdj
PiPsGMFKg2tyMUtAPArdVCCSk8Kjhsi2w44aDSleSG83fUuL1ok3x0AFAfkHA+8nzoBp1kbbyu0e
xIeBTiHFcesY+DENg3lkwlXh2dEWmE15PeBlLZy22/7O+rMQ2s5ItIIpH9V0BsCkP4EER25peHhA
rRoMKEA5LirjHzG9+mnhBGCNVbiROLxi/+bfkRA9cQPiOublM6ul1Mq5OBPPXlsJ/jfGyUIM/Qt5
+yIRix5fEO3opyrx9kQAFAANe5qUJ7nP9qg2E12k3lvkSfZLQ60yUuMksX/i2uaopwW/l7gqklUH
/C3TfPP5An3r37eWV2axGVo2xNQCNId8N6U5HJ8gd0qppTSkBWU1HCnYq2I4M6/9BmTfMMw3PGd+
0kH18HGmTGwys0sVU1Pslepilu5fn/UBjaOSjDONSHB8rpY3aoHk4pFee6yulKgpdfm65796EpKn
dXNx/uSFN5xbgjAAkroLWwQOzoJdNvytXhAwO8mt7AkJmrrWJ/Kx/jsY+YxSWKxqSbPMRexHZvvq
RGqbZU9OaE88Xf7hPTCmjaLPRO1q4uLGo4j0gwGZ/E46IfZ9zgiJpwBVDg8zb/3LT58nrMVjGMl9
jx9HgY3u4HP4i/iGyaDnUerG4mKc/2Q7po0Ef6PXuEkFGssGki5EVw0Wua+NsC7uLMGE8dPllsHC
rgk+icZb75w/AWHfYDhMoy4G4UPxfRKZgfbdXovvlYnDPb6ivq38Lau0JgQ1XeQsD5p5zG8YcB+v
a6ricvgFszS7tx3Br7PeNZp6ymR+Xc6SOlBXmISYnX4MKubUfLXQ/RGRgHA3eX2wtNlFcGW+x3hH
NTHFvy3IyJxF+YSoYCOrySEBSHckX94kYrTNvZ590EXFwdKDQSaYBSZ6+EkMfTyEa7fdNAkcp712
+4I5vzr6tCLMI4dHwWmSBYZaUcNSxw9VfZuUJV53R+aAdcqtTtgDKE6ODqtzSWMm15J96QgEToYW
9xycgS2j/heHDsyjjTmJAk7EZiSYcJOXvLpo5rdgl0pluGInQsI9/OBhOWnfoLGOu05vH+PQR9Ku
Kr8Nvjmgeg9ULRHlI2d8RMLliyQQb3lQItCLgxqzLNTJzJBVJ9Oluc8giCZYj0ZMEQ2B13qnv6ZS
J9YZkGv+a42svqOnVIqOASZ2CvE/T+NuCZJzH37UgzKAVmwyLNaYZdei9UzAUiSWe8WWAQ4cp7wZ
GbsEiHm9DmpwYsjhnf+gMpxmojETR48kVEV2eLlTYqlp3XpsvbObDuh7i3U85ShzXfgXNZFmmBHI
vv63fTS4p2hdNc1+zvfaQEsmVUDWLshj5s7LU0e+VgSNJpHAw0EDgYzeJmLKGMEjbJNshKLU5ojg
8Ola+PLyRJ4A2YPu0BIQ3UDyMFtfCit4gNR95vwO9uk/xUQ12nlsxnm6fLRnWTDmbBHYTWhMSqQa
Bv9jBbo5XaQ/il6vbA2MXnbktpirwamIWRldy2zRF5B24mEyfFRLChshidgqsJUtU77yd9jLe2sq
ezdRsgXhoPcdYZIfzvqwMk2hDokwAOwWE5DQcBilRnNAt/UQsxtRnigtLHtz5rH9VOyDY7WYuC6Q
2AP7mfxRS3/PqLsRw+Q+wteXNB2gLiyz1r/zT6nl7mjctnABhpIbvx2GfQQzzvP2KJUsYB577HYS
lfR4LUZGGlPfrpBXqz64PzjvAUSn51ZLVwr3sv6gBp7vqmhtNfk5VCf+4TnM2J/He52C9Rb7JWDR
+ZNPbch+G6fV6GIJc5niZ94cfZ4iFRZF8QPgT4HQBVaQ+ejfZU25I6GfgfNj6v6WUNdoByqWYjrd
Oefg+XYeaxo8HowoSu4SFiyUxsJFUiy5YP6JVA6rPbPPVIEspN6XiQnf6EKysl0o5VjJTl7VFxKJ
tBPp+sykYVhC7/f9RcQrJ429LVbw2N1R01867lxThariJcg3RXSwfzixz4rVjbGmLJPOZQtAZ8nI
uvAKzbzuMdfh16EqFYPrZ6/i6OZvMe0N6GmzYArQCR+rejS9rozKRJXq0bhuU4yry9lnmGnUQH3N
ktHTeBI4/VLfAlBelPeh9U7UsqmTz+w3g5ZOLLK7+BGEZQGNFsMr3AlJqfyw6Af6g45Nh+DwQW9+
SGEDQNe7kMdk/+XitNiM/AeT4jqUMsBaL790SKbhsgep0mKblGbpsxjd115W5AEiV+ilQxsn+t3p
c4SDVZsguMpDyVgt7q+2Si9kiIt6c7J3JlJuSYc3a3gTSBjrYTEQH8BWVcaFY2m/wsjFPuk7Zech
QJ5Tn4I8cxOsmBWFjxwRiw0VEX3QK6LdKcdXl3bCf/asNOLvd00Hlu4KxTBl3hmChu4UMFjaILIn
TXPN2tg2XFzSVI1xDWp+y+bepeUUctcjfgr+KjscNYWTOQOZzbDlA+SjhI438EL7wDYrJZv6cypp
lrr35dFf/9GQYL0adjIIMGq90f7NreWj9pkrlJPvC+PLbhv0pmMmNMmZNPZ8P5end+7oyMrqrtUP
1VDm1celJZOgQ/CabMVBFd+q4C8r0yJra0Hbx0UcRO2wDhvkciySJJ+ghjS5vS5/Hoymy0EpAOMl
ChFzt56VJdVskiD2N4D9cjGzS8Wkc8WzQW40eIV6I5sdDanzjoKdbvanPkk18yIx1XNDufeRqu/2
pcu2CqCBj47r3LT4z0hCHzrnneHSleeRpGgUycbZtZgBLnooMODkpO+YBSsHSdAj5UzMT9DzuTqS
PHRqkWjSPVnsUp7ANW9ws8Yac6EwR/jOhpSh6hUMBrc3Jk567ViyULkoyGjmEewiw/0xruKBxEuk
72B5rKCjlgxDcJMtU4tasC1YEUT0684jr/FGRVG/zelr/smEx8vzyyIeCdeK5WFwJrf3zFG69+Up
1w7NcJNllYb/JzCLWnCXDiBLPV+YV2OvWlqWogjeTin5mWAzBpUVsb22kqkkjQLeNZxYNF03MxlE
lerB7uYZe3akaAjlUgMrr4Dzf4FBol9VH/x5GllLBGCJxNnK5N4Z8RwUEdbI3y9qWjaxyRcVSgiG
Jgsvl5vQTVSYXldm85V45zNVZONLFVMXydjVMy0cfqGQwaCn+Q1bmfib+xkzUaA0y+f0j8Do4Dd5
p8P0UW/+eL0wSZX2DOCXN/2ORgEkaVXTWaBIK+KZxnhfjev+EEwed0apIQYdWsT/OjVlbfBMz0Ib
UeLhGoKYTPrxcf8tK2Hnz0FpZASgO6yxa6uUq/mDxpLwwrkPQST2wagAMEyFAD8aY7XAkQjAPlZv
vgcixOV23pHhRM3ZS8q0MjfckK9YT3ByiQXbFXdsQohw2alI2+IEJl9hkrs3JPzBKAA+70mhIyez
1QQT5AacxLSk6MX5r5a0Bhf/nNsNGzUsLRoceyybod3BwSS6Efw4nxFegrhu1IYkb2whgRFfua2P
J/329TzRCFz5O3YDkJM4XaiUJqbE0T4LohoF8JLYPBtmlWAMBhoA9kmaozwgP9vOzmihM9ELsy10
CK3M1Hhtf7gCr2/2gaB+oJdAjb3LnPq3uuhfwFBU8TPnao+MaJIU6EsOdN/38dvYYnLzdlu3LdNU
YndVbWQkXfQlSuDb4f2mGx/GuzeJ6xTeYUZf1G7P3PGgxVCc8Ipi9XPbvshPGWcRDZvcxWXalhiz
A7lo/AvJsSktjYVhdABB+/b7ahz820CzXieM1E9UEXgGysSUgm80/yTF+/C/9HF1iwIuWidIWj5Q
y5wB2APyZ22jblvVbIbT8QmW5oLP5zYAPvhTqAdvQfmv+jauD3goEHV7HRw5n9zz7Kw1d+pY236T
GV0v+bl1bBD/12kZ59KMifiumBEY3v6vE+q4T2OK61Kak9Wk0N8xWRCgwR+wyHU8LAT/hZbWJMyQ
nzj2duhoD0byCeMYsDkrYJB0pat0iPqBr8ekxquWEYPeXx4iRGWzM0KRIdEt25Oxa1nSeUjCJ0U3
8BTdMKUYsE3xY6ylCWmTiO1F0XhO9yGAWPkSDYf8sXdjO+Y9jUjwfB9523HPZwrib/4lcKCrM7Do
shYzQMVQonX/JQf0ZjcQXVUt0/P9TEJu7ulpRaIvTQfyWge/TYXOKLsw7oNXIVSL14wjbg3/RlHc
nXk6ZP00eoJc+VrKxhFtIsUa7q0Jl1SHmEo7YAIizVsT16ZxHgHn5asGc8qonXDCC3zs7OUOLhN2
zYls9Uew3CbnUCc0Kuj2OSPOEJNBEhx1odtsI3ttOKpnfeOE9304quXQfaBRmfizZYLGGsWOzJw4
Wa1mXQIcZ6wuOJi4yPN7XzECmtiRd//sFjguKqMk5nAfxKCrVkmDJnTWdqCP8omBUssff25dQ2Hu
IMPc4nmwMNXj8PCrACS3nY+x7Wpjl/F5ihMzQQwOIdDPynEXqiPcrQwPnjLheftnKQzFABHHUqQg
azQERBJRLD8J6tVDyO6fK/NuGg/YzI1MHaRHvcDdRwTXnOsyWAgpSPvdvC9ttyVaKuHH3W8KgjD+
GiZfj4FfX6cho0VcCs1ops6myNzfZwH5jnmW7VIZJviHca1rgRo05M+gemy1Z63xY1EPF5kBUbIj
u09W/7ugpEFXALxUJbq9kvUG6lfHUwoCRs98TDn8aPd2tEB3F7NYQiBX8MOhQw3TJOeXwrBiEaIx
sMTjtbBeotVmq6vVeZfUff2Nef7qxCvrAMCqho0ApvYIDjCoC9LzdWMZxavu0NiqlbNf0o8ddR5c
X3WRKR3TZNHukVr4/trSUs0pnGmlxC/2CIXSjv0NNhmGV2m3b1QVH7UdVDAEaNKcO7joqEGSRz22
KTHLGuU5mtz7GeESqoaOpyDaOf/W+bV+pPXua0X0JMG3V3x9eweBWMpGq0W5Uas0V9KvzVYbl4Br
wG9jkbU9Twi0079sOn6flqxese9LaPpPKoRAfdlESMFWz72B5Q2wP5jAuCc20mzF2MMrKidnLcgu
Ep2i40wU8qMldilxTKzhH5nZ7VOXIJN7C+KXPr1Ajv6+2OLGMKa0JSjEjzWOJx0W1oi6LkpaFpcm
qU8m0Tx9KwU/L5Y2EsfSJmTnjHXlPAh3+dgQ8ruQOFfg+u2TEy8x2UBnImovIMdYrGQE9I3tzLpo
jBnUBRpno6J6jFJ96gt8E4whlVjfFBgZ/EbOHSyf2Flgd9HEQv5OzDctd+JZ97EwBPj/4QSt//H4
RHhYSEMkXAJwigHEsufdQ11rHDH+LQgg6Qh4KtMLaB5f41mzwOL8hYKK7MAlkSD9xnz+MYltgpGi
hBpO5KWHWwOjCpGxE6oFJQUegN+B5Tzp/DiZVJm8pZTXOD0MIZBGdznE4E0ylIo2k8A0LVYiIdKc
O5YIv8lnwcBlwJZFfgc6tv8aMd+oJwAOEFPs2krdnGZ18jMcNga6ToDI7hKljli0AGjLsKqB7yg7
WqRPA2VYYxYSjYeBbqUOKHdQxEp+jR8YjAZdwHCcGHWZFYpQZyWgFeY2Gv1PXgqus5qc9pYRs/A0
6WFfO5uSgXJyglVpzsVdOgakNosyHgm3ZAgl9uX0UCVyVLXPIKcB8CmWND1Ifut8BTTo01fxeAA5
nJ/5fO9dfbKfK4y5Lptm5hM2MBVKl3Vilx464e1BeEEeSoa1+GLiIITMjoLvge0gMRK8ixeoudU9
ppKVyzDp4h8Fxh/F6F65Rni0l8vGB/DuB9hgJ2gslBvnz4e3XOX/yPij14OV4f9adskst+gT4rMO
eA1BcSWiXusmbqsX3g8Z8fRD5TyzJTNKkCcB1TEqh2lbQLsfwg5VByHr1xtsPRd7ULLBTeyLF8TT
ArYVwvn4qDTXwycVx+O4IMrzUooE5BklBnBgB75/EWWoVvJQDdcLCkrwW264/zODSKdDf/mnJ6Cy
+vgbfZ5evCxrdiMP6wt8zexnCQBlv0ihz87oYjnF8Isbsva1jTztd9AwcuFr4W3gFsk7pjgyfi4J
7fWopbaH855vpq4Jxu0xUUdoqLW9lKm8oPATJ6tpzvkXxpwzZn4GW9/fP3RMkIN5uPo9d5C3VvYG
b9OENnRBhd53GUTjDFXR7EVO7QfJC0A0XUJ6uIs4tj1osanq7SYflIknjkqQCbeFkz60RHSrUm/q
Ckz7dAIibE7PKA/yPqQMKEUXpS/7AfolJ9+8k113Jsr4Ui9gHP/3+CWBgD8H2GmGetITnEUdKXNI
m9rsekmeYk+TcJDaCzObcHVYgyNuj94bRI/zSQC2niNNANG57s4lriI1vjAs2Q5QREpz3PdHGqNg
N8G/wIYWevap7fnmimjv5t9QMmfEOwEMjnUT41VFuCrEGUa+K6cI0yv9p3wRcSZoGYDRtaHiNsPr
y0OA4P7RIm7ibDqpMQ8Rw9y0ofOf78W7cE4FuJCjb3CNZ6PqM/Dd34yocSr3b5jXOqoCZEhtydXQ
s3eNSA4qNMC33d9kWdLHrhnaFMWwE1RrzaiAif6wt/SsBJvCeOtlodYg79RCTxvwKSNpo08c/r02
yjoveM+5QYSNotdaE+M07x5xjqNENpVva/TaTEpR3oufqxEN/OOTFffMNTAtkJs9ArD/v2Zc8QGQ
qyraY1zUXnQjScCptyB1Z/pY8kPIUmJ5Q+Cb4FZ+c9xgcQB4Fq5aGeEVNQDIKcX3mcb2KkeIHuDX
TMfGUwZ8rytj4wnSnffOexOsb4ZUJVNeX4LJZpNhajbs7tyGkya0uhLsrVJLkD4mSQRtJQL7BADs
Fx4q1VU9OgQjoVqQYC32V4xQZRwl7S0mVfYi7rj0/Ef6xHkkoSa0m++rTeRqCCrRWyNtHb9P0m3D
pP27ssOGQUG07foaDOqSXbaLVdu0y6Tnl9zCHKyUOCq/lhtmJ82dqPN0ZXk4doSYPoWNIywzB99+
7gDHz9fKAHvB7RcutC3oBqbdlx4FVFDOB+9c4dThiuAu2BE6NzddMmfL68If/1x5e/Lb5CqOY+QW
EbDkd4gL6eUtHW0/uYhHxNzXkRX2jwl3LbWuwyZmliX7d225OkvHD4kf7y0HrN1IHhRMTTvLbE0M
fydkNvbcBDEEjEDueMyI9GIK2js5KOly2P9sdB3mrqHb8L/yzHaYqfLOE5cjGKTCG5jfR4KQ0+mh
gVEDz9jhKhyANasjl/w2jhbk6jNC4k/bWl2GbYhsSX6c8yL4naku3/4+CjNExq5CRxL4il78JojM
gpgMv9XrQL6/SEuRm/Ep4A/RwZkpCXHbBfd1+U0Rg18JBAuSGRNWSa5ycZyYvs3GqXTDEy3FfZlh
GzUi77b4GX9/ajmpx7rhjlVGWNG83B0iz/zA6jFTh7jT4yWwnDO702F7BBW+CYR9iY9tFHxL6gk1
OrS5MvC/0Yt3pNABE8esrRRvttRINFyatr0R8L5/0Y8xyp24TUeVaozcTDJ3kwlpq7qaoZXoxyTD
sNuq11WTjpsZjZF7Uk7Ze3zd9BMseNEwGjAaIXC6zloaMItymE+TdZ8els1qkEwynQ0VmirvtpOm
1DvCAhSucoTKEkWuhhlGEeI1Ge2wer/dZCN+RcKKXzmon97PbfenSXdBYh93HfqrF0BPnx6EcJst
LMroLIp0iKc3mWLzbh4eBUrKTCBrwynZNMEPS6/PgDqJrlksjUssGgDFBQAndfkTHiE4pbf55zMF
QG65UwOsf+Jb1N1fSZOSFcTZKWvOpihnFq5/uc1gq1quxG973ET86i3emhWgoHmNt3H/u52hwT8P
i5TzFxJeUmFQpd43cA/AtHbh/GrBOa7Ll/nUaCEvkZ4MZcT10vs4uJHTttbhTYIXYXArJwEx/L0u
fkjTyv0Jsp96XPqaeYyTnfb9IL/tVeR0CaWXFZnmYG4GCICcaH2KHvZd3tGYoubhA5jS7fM7p3Fj
IG/LHCvcnnYZV2WF361pJhvHYhbbaaihWroD8YKBuJY2VXUA9ChkNuUWOzYhO2mhVfGLNDHdti7v
R0rtiCapdxoLZKzmAnwV5Mnd5dJjkml3XLs7EWO5A+VvcC58VQPd5uBsnWc1p42R53ILA8BpGJGu
Pc3XAk19T7g+KNijZz56O5iow/xDZrqeIZx1wdcvY7jrxqZd/V8fO71akwG1++WHucnqeo3G+/qI
Ul/FMZqMkN9SN46vw4stN0BRlXTTFMfa1mcXvVR5AOHiqeKzGPm3IP8Ti6Luger+gDHsqpSnockI
fR4svge6T0g8KBifrAy5U+kt3Ay4sVECz2qIvpC3P/EGJ8RK6j+OW+XjRTsVu0HBev9qk43GuPMk
RBGTF012N/KbJmwi9nce/i5KNqzLY/4HuKm11p7rTRe1C3/6cOU9CmofVNv5YGcstxC3xiv0FZ83
gjT7IqfoCCQ7amIQ3WJgLOT5yglw4vvqvNJ+aF1hd9RoIGi7ZReuwHBZJmXkpBznHAEV9zX7EjPA
S9fYqJE1slwdTCvo6B787nsptPVQqJjUmFVWhm9bQAj64GmsSRofkpqm/eMslKm384lx8aYs2V24
e9tLF7RIkHQEr8L1bqQHIptIrQrW+Tz2JZIb4oragLKx+0xDUK0Xkc4s4lPEj6BJyOaagz3wPU5E
g0RynLFZoxnseF9WG5fPETNnOiDqZxbIhrdz84Rsfk5s0NUy2oRmclLUmsh4gcYa0tx4vx32tNT0
pVj5asdFyE6BsnwiqGwvOn/eLUDHEGx4rnZsnwr8vf87404hpmbE+7noWuUnAD/BDjSqpV6RDkLj
B8i0vHDWff9qwcOUEAlsHmwmkjZb217cQHqS78kJmIxtSm3xBeDotPmKgDrwqVokz7elczkT8DEq
rqYw0GdG482so7VplCWIRwyFb5IMiA8KM4egTOCTtQ7RNfRznB8cYhJB4sj8qnXH3fKvRHVu7ZQU
n8RnJZSAw0uZcksUMeVyK0FdNU9F8tuTDeA6boI3ANCufm09sAK0Ns0oAi9HnbPs/AWXbJytAKQ4
3yqrLm9PysDhTVIOTC9Vg5PR7qEhoqeIpKqnUMxjFf4QHCY/ThEhm8d+QGUop0dd8wz3bc8Tr8vP
kWxROeIZJNshkPu2M1JnGFkI2o93W1HMHJc0CjEL2ePA9SHLWVHp2DSnAqD4+a+ZZFpma7ZGsu7Q
VvzWzUPsq+F19AmcY9VRNA3X3LuHyWPAM9GNJrJQOEWO2YeKCT9Vw9pl5taZpm6DBIYJ5Rd2rqIx
Lgzi+d+Bpt0h6v6WDNOS8zTxYl2z/ATNFkRbek9v76Brn8HALZyUoYsw4PFTxvZxycn6XPd5uUx2
GTulGISoVgN3asHE1NfuouLAztH2GTAugowcxAu9E8X/9raVeLwcZbpcvMgSeQhwyNfoLQA6jLNM
6HlqAgjdABfEmYV7C3Fr8KxXH8TMSmSg6Bq+hmMQtSLNgg2fZnhukQKJmJNW0ZAzRaP8rvdewHWj
Dz5lwkDq/MsfhGf7oXP6EiDRe1sGJPS90GDIoLeQFtyKw6ykaQXJxaN2kYTDUsB7YdKcstAkeXf+
IqskjGbbfFekRUzp1UCSQ2sS9M8MKnSiKWVSut0w42y6ffrOtxrLtuJrJAhJMOSy7IgAMpZGpHLM
/3wxg9cdf52SRspYZlSN1ep9N2vivEMzBjhGBXRfJDyQkQyTSpDHh9sbw+RrtR2T25a+NaiKDuiZ
8cW+vqKPZuMUYJY0X7G92A9j+yBRyh5U1V68smWsYrBpHokGFCFne+sWgEpI0vujs6JD7i/9sBiZ
yGyMMV2+KLTD1Jxcy3BaJZ5YKqYOOTAimQvl+dT4vpmMs0Bj1bliQ/Itnx4vJ/jlTVLE+RH41HIn
65nH9ApbJ9iQJIJluAQ+Jb3TAg2arhMWICK+9ZgOFAX44ST9s1ZAf9vw8JfWA6OoN9luxRjzSKeg
TA+ZdQhISafbFdHN/C4kYNqWWL6c6YiO0f53arDiCz2B4s66ccTzyJFS3EFuBcuTQCkfuAORRdhD
r96dqsXSOasS3U4BNg0/QmyzJxURQFDBW/A2lR9DvBwnA8la8GKqlPYUa3UgZwOlQqz6rd+hhDVP
VY3noXxUjwGiBXJJvwjppzHfDqC18c/b3I0RERaWe6sEd9lf0zaH536kCe2+qgFLKj2afnzDL9xJ
c8kNprHdwnlF4dt01F5LoODvRXEwPOO5ZZ9kNeQ4lP8mgkcx5fIXYyUPSfX16GwnrT2ODCJHyaqX
YmmlhzKAeJ9ZlGPovmFFwZ4fFZLFGwoDvUCrpqTAjtCxRjo7XsFWd28C4xXCM1DkpQwR2ZIcjkF5
acbA6+OFvYA4tXcuqZWJC0LLSNzXVGaXJKWXGhPrESFpem5B2vjJ7ewF+TZrlJwlqCNJstyg2B8r
yP9Qxh6XVfqzOfYNFbbUTRhIzRZfR7KrW4J68KkPVgHvIBfyBPXZCGfQKMR98UnNkNH/VWhrAFUQ
XR8mDkdOjFPm0ZaWI9rgF5aVhFOezFZw2hS3igESxW1NitBdgJdL76Lro1mLn4zuqlzi9xl8c9yf
e8YoeipcOc1iEzp3B+mapg3cWzvwPn0AI5bW4yWQqbpi12XeqoztB6enP9q4qolRQC9kC5CGz7gH
LdX0rPU81iVA/dvej/4y/d9k876aoAdPjY3ymUCI/BBz5VNAwRZimOYRgb9O+U0X9x0rYge7th3j
FX7ykgfjLc9/3cPyFdWstsI1bmJ/yPiqF2c0LbAGoCEfIrAoBlUl3PUmhsX8muJAKwIV9J7y0Ab/
JOgf3GI5vsDdndCxgPpJfu7MQn0g6cNKVtkDiUGzaoljun0mZI3Tq3lM9oiMRcDoQdBvIG6I4CL8
o/7/yHqAcBdf7yQr3pLGICu40/nA/epCvhi4LHtm5HpF8bhVpwzUJz2ioayHyDb3aVIlOTC75aBM
oIwwgVEuh/tFKakhJ0vYNMAyqHmnBIMQOdQr+DCOgiBGG1mA//VrFxa2Yz2PCL0oJ6ac/FKzOF1z
DFN5mhlqUAZ/EMGvBTqAUutwwa87HfsKDIxJb0vGCLH6oVRa002pwiLyMqcWiSIIc6WzSC2uMo80
TDq5UmuXfdZoNnFESSItlIxxbMZKplxpZx9QVCsKEm/WsEYEHd9jQyCBvGe3tte8aLCa1nh+31Wz
GV9QrPsqhGJJEbmupj/kcczT/xBiPd2NuBZOPdjUHl0aMJYXYnN6e8vmwqInq26l9F8Zcx10KSHm
q6tU4BnEIZ9fZfToEqNgXmysPyaKnty0XIkgrhFpo1XrQzYAnfuYyMO/eJa5OHYRIq9tkFGx3p3w
tFEJ4O4MM7KlUaPn2gLYby1vuKDqcIScYje8Tfh30RYua9UzcBgS0amYVd4ZxWnChDv4KEZJ4wzN
NvrvggChrd0J0tHnyVAzPeQQ8WCGFVuhIzjQUxq+nqytWj9VAyEnCyic2QzktozrN95+C3shTqR5
BmJ7V2bV0a5/guq4MUWHGG6+dpBKheEDxaYykunK/Je/xsQ1a0/tNuIwdubN1Z/dVLey4eRx6Qj0
X9H7V0qX+q4XQMX+Bd6nQycNYO6hm1ufq4wZFq8vxLoYwO5HAcliIy6lKqWIEpJtoIfMOjtsovQp
yqJzAf689WWXoZvNb4Zye+EsyuqFNeI72tDPJ3qXfSnQeCmweVxa+xposW3qUZCriSgVQN6507XX
H6jYhNWomuj7ItSbGihe3PsypRMGDU7U4jD4/vQKHjk00PjGrmoRE9kfLuXXbmtcWG/06PiAqnf3
eUYKkLzpmt61PUchqAIn6Gzpm7X1nvajpMvlD8USvqqAKvRgyUSjB0B3GZ/TBMn7/a3HFE5XIksC
2VSiIL4+SP0o/I811BgbwrBLIKJuo8wiPnrTFWk7iqjRoiM2xy0UtMjA85UmqBjrzOWbRGoeEmFw
cyyaYVSC8NsUFAgz/h0d9XLBRatKQ/HoMpdjsI2uDZDCD9zbI+EpnaIY6TAU1NgFW58fFGQ2tIMv
coPfByvjhaR1+J+iOUNQslwhn1+POanDGGX1jhpqlC7TMxpXOK3ytC1I7P7IeXW6nX28JjydFS7/
aDU7Gqr+YU1ezh848IrxrQy90ASEptTMuT7ivs3pddA3nPPsZfeofptbg2jsnYEaXD2AlfVR4pfc
QKTLob8R3o6JZYsFVP5F1/0refJ2O41lVxgWtyb4JFYMbG6e7ut0bmNb2oj6f2PGG4YN0mWIbXNK
fnMy/nWq2vrlrkOko5yuJ7x1MGoa5iEMCo/0hEtHWTmB/R9OInRPU0CUUZ74Ut8IsFWcUFOr4Xmz
vrqXuQEIOQ79N7aKAB/lQpB351PO7EvPmJGDPRwIQjmGoXkGnSEuzLGoLHVqXuo+9SFU9F0FtrK/
4zs1TV+WCUAgNRqIBfuunQlTSu+8FQhG65wd0/cXEz3MkeA4ZrBTEudiB30OGFJxL/+SApUE3hGo
C0uw5PJd0IAr3pTb3TqxQ9/PLGgscvlC+vGQcfm4Uo5yrRWLyd2Tex3XdsC/+UWjJjUDC4qIFBTP
wLwpxdC5iT/VIvu8fai2lLUjTVPW+8GrV5kFxCU3YxZOhHUqQS2JcFpaPVoTczYwQF2B/2FC8yLK
iX4tLhN0kRb0f5ciItzFulSaLHV8Dd/20x7AvoAbI3iveFlCnmfuhoSKLry7pZkHrvCKxvqf108o
B8P6JwScVWfeF9SlJpBDQfCmglfw1uVKvei4Z0lVHknqT5fGobBOFWu6J+c+yXSIJbP3kXGM+UXf
FwteUdNqMusEi1pBjPT/586bOfcs+V6B3mK3LhMIse+PeNp6cKYKhHbXXqC7ODSFiLu/yhyqKMqZ
+RbttibGu7sQbCaPqDXl/RHkwKQAmk7S0LDUHMEcQRphKMN9WWWvPOZjE7Z4IkkvnrALqhThPilF
v8raJX/u1yYXkH3hhN7Ip78b1f7QhZR8NnHYQhkOlDIPUhUDQedhW5uPP6af2omUtf49Xor5Sm5Q
UwE2e7j9UHj+Y+BdiutnOSA3ns3dUQ7rwg7AcyJsenRduKX2ge7fIV3ybfQzP3Az5DvCDe5NuREE
KsyNCF0sQdDe7RvEZVfkayk9tWuLJeKUBDDu/h+xA7OQd6+EUqRyKKRM+GWQ5mF0xkHvLZcTJFHT
wB5Fh8FIgVei7jytbNeTu4VLHALmmzH4O325aTyrA5QAshXmg+ZI74I2FHqpH3B1BPUaQfNGHEzj
aPyK00p38HGIcg+07Gl5n4wK64HHN0UtHdTQ8grzhQNTpny6CIKRNvHK69Rpy4wE8ZfA+CcnWzVJ
hS8xuQUwGRdRyNxv1isEUANTzUSwXI/voc9pu1hgfXPu0EDJEH4zZBcwd7NpYHfXPgvlyijBeRuY
iTJOA2Ik6SjNK272VNyOotUMWXZnnOLMZH0/3Nb2HvY2WQYIwNRu5TXG+BU6jWFq1gbZbj3nr7AW
Uu77aM6NfqRlhuiySZYJYm8qgv2nT6TzUK5Z1ewhrv0suvvlg0Lq/LhIKBCYIlHWzhBrkiRIzxPi
xetxsYbv72xzwf4nzd29XrlrwTE0pjSYqrF8cVwJCtISzLnVpJYg0fSaU7HoW+4voV/OLNxCla+b
6XdoPDbC6DPCmZFaDOn2OrofRPanA6WvYCo0+Yyq6uJQuZD10tQ9WmIfXb1Hzlr/mciYriPuOnZe
53vT5HaAoOpBa/7gc8xPerb/hWh47gLN9D28YGUajeS8AsQHqsOL1f7dLAOmYsgNCypq9eUyF4dn
JtKJM+1M5bkNBFUyb6sIpzT1XAqb/5t6iAMKEAn5otj4MlK5xgd/K3hMCw/DgUMk44KeIEy+Sflu
p40t/u7v+eICMWdCwX2cyPY9c84C2Nsxncm1zsaqF/jb4/v6XnopslT1JAN0qVtOuPKgIzhFdrt5
QBj9zlNGPADhYCUe2m5sCU15nHNgxy217FVOgd8/suCub5iBS7wEl9pyIJMayHtSbr03BeUZyq0m
6o47k7kF5qzyIIRJyB+xfgMcjvTOCdpedFhQsvArxg/sNsIZUDLeYrHldUNdiw/KVlTLp+hlRQXQ
awbjAUfjY3EZ5YcJe6rCgpKeMHYv2ZpQoiUYxsAZSsUG8tSlIwG9URHM1aqC+nrQFF+qmmXbSJis
vRRnF1xkBjUlBklPNwJs7O1yofR3u9iww+wgjb0sF2JyZtJbjntfLkCt1KSizXFYqLz4YjKhCw4D
bwTWGXxiWZwU1TzoVW/LjydATYfr+Htm6HG9ZFmEzXoTTo65qNAgWC09FRUv8QM0+lhz48Jdx530
lS1uQ76HSGJCbHFWiNAbWTKzvgTXx6B42fWOUxDPtCH5Gqw/TdiyP0xulQGd6St5ssIuOryPCNj9
hp6r0eT3u+KxyKybtxkvqYyjgTZUFfjEHvMRp//b48T65/RSEtRLurUtijQuhZncOonoj5IO94iV
SnnpXLh+huCpOoQ4NJz3UtgqBEPTRCzo396MZ9yji3J80iDgAx8XeXnI7iQBJGiQYOQt4xZqS0iI
fsjxBR8xUZtpo42GyjStXuEzziPB8sJZd5M8kdod3fa4IAcD2VTr4FcGZI+19gIUvH2k+wRNfJxp
ehLzaeVSl2uD5Jyy2qZJGcss3xI37XFqx2PnC1me3E5H2EubnHpxtQiEVSfJMvqrDG6YMEIfWOrP
+CpM9q2yoykCbOz3MvStheB1g1ZpLfs4cOiys6h3+vN2o1lHsApVqSfJJkRth+k2Nqv1VnD94vXV
9jte+/RYhREYNgpsko0aQf6QwoJ8ScS8n6VbLNTYW5JROTz5Ql5V+xcEraCptdYdDSM0i0M53mP9
16qGHo2TZkLtqj6mnQ8W7tPKP3G0rDTe7nkVQvXaYOqzyBR/MIPZ+cpaWeFC+AhGbRxhuyBk2wc8
momotIj7LSoHOFnpN68QMdFL9p6n6fOTCXS8UsxpPzlmJDXKDbQjwQE3fZDXslDi6fWYpXDBrlnw
uQ0gMC+s4XX0XIvbfo73Ek91Tx6MnuTn+3zh9oh0Flc5MTcOFKeqfK4K7IUi7ySQGtxtWtUMxPKB
BTvzrb0oi9QRNjUVXW/RxwnB1AvR47OVrnEjp9YjWcdhXLmBNZbiGMAjaxjwjhS7BX9ZJxJXr7jE
u09sKvsN0W+ICT7grg5NST/oeZ3lCpjoTgg1EouJPTqbc2Qp32/6ptSDI301JKFkA1FIxBkR3dtq
F8auHFEocoK4MLJo+QHpvdewmcds2HEhnzcd0HTS9MbA7uf1+0+yQ/XtjAPwo6y6QSt2C8cD99LP
Geczod99uyZdxpLvUs23cR9N5olGDeU1elXTFnksiuGbDjOGF3x17VKRFkZtr9wBzHlGozRvPSWm
E1yWFxDFBkQ6GC9ZUpk6pXwDenvQhxdIKtrhH7/osqXn0N37zUf/jlSbECvuCK+eDRFCuOticG9G
8M0poB2Jpy6nLRtX5R+mQ1lRk1h6j/9UvBXkYl1sWmaDEHKPBWGj1Ds8mgXC1GP8q9RYvG+7c5oR
nvgA3VrZByUI5+pTye4om8qsNrpVUQTiNGYtiBjEjojxPJsg654tYio7no2qz5BGU9UBuv0eGECQ
gwGtIehjEneULWOA6Ao/F+NLsFk9L2DAE1lohW7ZljBhE4xuXuWH3vk01dPn/YA/8N1bv0WmTEH+
f/VUSbPoabcRAN7w2itO+4ned08NGjHNZ7bsgYYOQx/SX4mFi/u/OgtZObEEDoMLBHN2O0GWTRUF
fHMc4DQlgpm+DkvEOyNmasy6waQ8KYI3+ka1EziDt7wRta/DXe7Md0pVTRVcJQC6UwDKB51fBpb2
Agn+o8eHrHhuca6cxWnsVtn1ApBe3e1qMb3CfrRFLXQkHSFSiPoiF0mbpp+lcokihAp8Q0lxvIcI
T1+YbDZNkpMaEW1zms03TOvt03cc6C0MYqqGydHXlGXvkzGkPWK+0GL4CNpW0YwmtKZZWF4/yWQR
IfygD23tjNjGPjZyC+yoq/AXprawDO3alveDWhjbjPU3tbOebG5iSHd9moOnc/3O4R1fc13cxrzn
xyBtwJADh3aSVqussxWTceJaOFHADohCH5+ey0/jKcndvm3j4/+Ig18j0IeLdS37P5ixTWNYoBjO
MS1h0mPZeO8LJMcPZw4tXzBfc4hherJ9LUpQ2zQu1q8Co+6JTatucj3QaSolwCNQ66fhpMMwfZrf
SiCd+imOomA+ydhQcK/e08vGpatV5GuWTk1ddMzrb6DfYe10zo+ajFkUYQJP1uv9Y7S3bTuxDrGM
RsxP1Zob8xU1k5dqathEGh2/93w6wEoYUWBS9038JJLsa4jdZ8Faf8e0IoqVMDTEz/ZK2J0jPrzW
vv51HH/9vvmW7OCK7rDpVjPvTToFJNbNN6vBDQF9KfG961uCCPA9TCM39izs+GK7DgEuRY10lssx
HUOwvmzslhAtSYVOO9Fmqk0FF/ZzVqQr8iKz925nwYmX1h8KA7N768QrgirCzoNU9/93gN+ADQw0
XL0JGRvA25CfLb3efm7gVBflPNXsb2yn41ed58WCyQU3hki6bcFiUPUxHfMwU3zHroMJBESTXRJE
NiBI/GdqDkuWGk2KHQao/tZ1DukWCUNOPfadZeVE6NNB7F8w0RlRgz9vJ9GVOq1+8OiE4V9oN1b5
O6gqxjqFXbapti5/4BucP+RdYSeIAyCo8jNONhNXBOAUXySjuaGfw3R4ELe+s+KOarznici4A+Ln
lUI/8B8sO4c3tP0wgzZ1rXdljyl7+gsEYoN9VqU89Nvgb6aVbvppe9uiR2fSPd0YsMUdkKUZ4jnu
ndZLqgpyev+fOhocR1ViQl3ZI5t4yPLGuuJRSaeX6aVTma/tX1tWhGRN6TTuA973rIS7ERhbRXei
9puE0X3Z+h0uoEtjl11M/6nmNV7BKm9wvJvxtc+uVVbn0B9xnJs8kNGLCvzzCcn2EJUYIbWJ06dl
onpxVkfb4/X8Bjw5mi3vlZ3LrhLkzmODUummn/7MLn2wZCmRh8b4pdVyu41kWRY6BcUppxnEce93
QVZobCIUCnvWXR3GH5OXc+rADlGbDy4p+RKVKNMJbGfWAyrcyqtDCZD4ejgrEYqj/BW0OAkN0S2J
L5ALJ5R9gAIT42pwYXJh13tad9cz6u1Kcgh79QrnyqsdC0UTj3TRtW9gPIT5g3spH9hK46gPF9Fa
PxVmRPN5jczuioDeaADNk0EcStXv/C0V6SsJxkgxjVYxk9VRRc7sp8IoimuiDyeUG4+JwsdGn4ZH
cI7m3F6qcDREDAi4o3btWFW1YiTJ2FuE7R0d6RKtR7k75pU5V6Rm3X9U86uBgx7Bxf2U3/k5Ds44
jLISVmffVQOfG7ipyn1JtSEc3CmFu8o79nM7p6Wv0eYov5J0qMKSIOHYgajOsfk1Y7lAB0kpXxGQ
IZxd57rzJrt0ri2hEpqtJw+Wc7HUvaZgkPHnad1EbkaTbS2zW8tLtADWCeowYE2B68WZTzEO+OD/
jS+Hj2lXa3aiZaj2ZAuSCgb1wOf2gZJxHxIKe/T2dE2b9yasT2WMntYbpJQ6pK2+72KVXcpKeqrh
bZClsB2z5f9/plBSl+z1T7yzU9EyvfIreBWqt5xuF2L08E3UQ7rSeu+8Rg3YdJ4DQMNhYXUDEypx
nYqUBLolYP5Mtvx0o5pDT4mlwCIsMzKnsjsP6T/ev3TclmkXcg6Q4wF7ItpIbu+JJkRq0eXkslJk
VNLORjzKusTQKvenPilVpwVZII2wcIQu2Rh5d4khQwHraPt4rlf/Nxxd/m0nQRyl3Oh1ukYEgljb
CCupOFlWI29p1d4vR7EWH9fuuSrNbj5NSgQzcG2GIhINu3NLBIhL9HjOpp+m8Z1JHID+VRUK5GJU
KUgY9OFV03hquUwOPaQr/0K3aT+kixIkByzxAflah/Tb8cG522zpgb5ZCYhbFyFPhKy9BONBcTiK
BmPMsEYLWbVPlXCnKuRRtXcYdnvtwJAeOKwXDhjiNPYK2K9uvw8Xw/ktZ+Ith9EED22Fy2dyuI9x
iolKskES8usOZVesWO5WLW6SauoG4ZzWrTO81O/spvnD7blzz3SfTE7qychWVuz/2Qat+BrN09ts
P3vjGqySJqwM4xtsJhvk0utXlu0dC21Vkq0W/bM29pqU5k6HnBiNEWka9nj+amvcbeNvYF73HiJz
JQ7ZudmL3UeoFm4b3RHpGQGiF2HH/mGHNrl5Trk70dfxxxFF50Ji/oR0UBawjZV+vV55QEcjDdAM
ZNq6F39K+eXqV+c3FjvW64ET3GizoIN4ngGjCjvtElTQXiOJ41RbTJ5vO8dUXaXYNAbsyR0QwnL2
2sW6LRnyFEbot/MY5WtFuABbccFhPFYcYsBZLWdYThwqOssMKjMApcmdVrpppWRCXDPzsxqD7CQp
VvH1Cq0hWBgRwJgN02mxQd5xDdIUD7wMECm9KzxQ64eTyGJceJh1jS/FyvOEU1Lz4NvYmYmqGjix
MdmSk2ivQPpMcTIkCjTqCSLGXekGe7DNRDR8YqxhigkhgC2ZRUofmoONRzjSiWQl7q2xyEXn4QJL
kHmIU+i8nI8RYgErZ84AQNrm2FAA2zLfxvGne/CJ2M73zF/Lg8jV0xaLhpJFk2Yenh6L2+ImHwbF
xHHikU0rW1gWpo0/BvfjWMxvzML6Qpzey6kJPmdtcvGWT3Dm+i1Km7DzM0THhfMHC5gtS9ay7jUb
wsEy+onr1eN8UE3mAhKkyMDsVfzpogVCZkvDwsVocxPGn99ha8+DDfpPpHnPww3WHoivlvSCMFoi
y6gzkdZ6HN0xSIw+ENCdhnVL7epv7TwC4xUamVg3TYADgctzEvVEqD+h/05TpyWLbcOvzAQdQWIr
zUAmfBIiRAK9L/+5sXoFs06DKSXB8sGaYX7mpHEZSBgoQ+dTKXlv45l3fr9F774CiwHD6+fWWPel
YIDrowDQ/MgScC4FGUF8w5N/OTcMPvi3d88d6lcRMueGWh/LVdDt0o/OkGcIXY5YocJGA3WWn6r4
HMWu1dWfw/k6HPvy+6XC6Wz7BZzk1rGCsX2p2TLDvzFuuBImwtvjc6FUYWzb5ADfMvkezetSgkj5
2s6BQT/F+I03n11PpPC94Z+BlG6Ifg2yeP1zdV5tcPGkZp4W4k2IzJiyxAfb7ACo54zaRnk9gXE+
wKvvmaKIbGas+Yx5b/HKZE9qci4HvT68zbUya2rV+5iCMLJaJxcPF+ccnUxx20vfXzcETdxs6Awm
9J2wVerUv+Y2EfWI5thryjTzg3chEoIEvjxRNYhWyI9QhCNGtYbvha3cf/OyNt1jR/31duQYPkjU
h7r86F6vyM+E5cordmoyyBt7Hwe7wmXTW7tZjvcrDlzqZRv48Hb7njSpSDXsoooebopeRQLqDNzD
hORXQVOXqZ4j/eq6OKHHT7IAtYXp6KA6iD3SCOCFGLGGm2g+pPiphj9rsyO4qxlp1l5lhxz48tDK
RvDckagVj041IUgdOarFmrFrWyb0Q75XFhyhaTDuQ0QHaSxb4HRAugkAqY3E0T9gXIypV/kXYaVi
mChBzSPozvcHMyfrzZ1AvJ0GDNlw0X7BobNtDK6elUFKZzhzyD72R37a0AuAr2D75qPT/NgX5dpY
EQDTdpaHIJR7TtabuCyb3np4MYuG/s2wCb4429gVmEol4Bkd09fECEN0FufCBFxfr1EjkAxrOej0
/Uc/z3rQU7D8+JXcmf7PiIXW0TbKywMywClwmyf4PGnAEi4novgCtpY/5rf8TOBBMccGMFbC2ZBV
ZEvoiuucPsiZveUBqUivfKMsaa2ourI2WCyvG3T4Lk0yAskoeidmGouLiMioUJJGVIXxAQanvzSr
xoK9TPLIJ0HHCxGebyKUiZSsZosv1gCQUqMrS391SjM/etuHus/hJaDQpCiDmJ72RH/Z5F0PMqe8
LAvMJx0qkqw7JmxEqDSm0xZ+jQnrMsCwZYfgFQssyovtXIs8nQHX88W3XHgQ/son2aXzCsSAmF52
WPeoRxZRUBlbP0hNPiFfMLn6d4KJVYdENld3xKRbIu9lvT5XssCiQ+MwaOB+wQLxt3BxuJl7n57p
1QH/NZMPAd4Y8kVPzyWx78nJRKt62IP2XQ0tMYa6bGebmxA4om98C6e3t3J37iDWjPxMohG116em
4dW4JbuUIHaoGtoLsRUqWo8eOW9tm4RuaJ8QJg801TUSVbhdqA49r47UQfL6wh2jMppqh9CFTdbR
t0+gmNRoVN0Tsp2zYN9fYuyel7/GZ01qmz+jBk3eELwJIbU1f96OvHH/y6mor7/abjKSeDIMEm3E
Vc9Hspw451ZljArX2s3wKu5wD8MWfD+A8J5lcjHROaLx57qP8BfXWohkUgJrXbaEX4vXASH4inYb
c3YBVcnNMoiuguNEBQfpWA4RuTWgok5zPYfa18cBox/KzNYm6yfalCCSZT0T8V/CCKuYE1+Ba3xO
7QtKrDz/+ddgMy8xbArBdn6kCs1sy7rsCY6pNdi7rkq8m09OhXehHAi6ZUJU4pB+WPRxjVzXN2Yh
mmj4c7uCfK6Tj3n0vQ1CIHCIsFgBhr/VXeljQYZA12FC4LooX9NbuJZWgsz+U4+2jHM0oR5qvzFe
m5LLsoWMrOajfJviNXjXQPljBuxbJMZMdnSJwsF4GVbzlHrQjwUg6Aa2yIGmt1FBDtQP48abTm7K
HedfvSojXlC9PLLsJk3hyo5+7MyGDRHGsK2zAkZ/RYJaksEVags8fAIc8U/MvlKlTsg3l6HKdnT2
PNj6ADnGKeGNxq9Q+IfpRCy6lAWReG58KGeiGYnnVcHQxgMzOnwfE9JJsmIPrUefRaaPVU4qAfKU
a7jbEBmvv9uu9/M8GD5NUK/DHV7Koo9nle27YClAh2yR41My8OkOXP2lUkaT7IGeH92TOcaac1MT
I6V7Ck/+WGiMFDnB/qNceOGmRQDvN73eZCu+ivrRatxOLfJc6WmbppHqykId8n+ZskF/a9SprEar
tBLC8Iu2LyU/PrxUrbldLhGQHwjT+aD6YTndaATahd27iS3kIqk00SaX4Cipi0rHbLHkDn2XWQbl
p51Y6VxmVrN5TFIJ/VLalwUehVfd55CsYbxgs/AfxfBezJc8GzpQDq9cbSN/1C7EJft+mW1zEXoe
5iWWJdT0Rz3g6rSh8Dy+CUPHHIec0pBBWfKunczdkbsyIDNR+iYD1DhZ4CNH8yW3cg4nRJcjeoLq
qpd9Fp9qqLZ8W6WRbJeN250vnWVS5lhdYLOcM8Jv55xZGpJbdfjaCS6XNSqf/qemMQJXBU2noZJA
lxQzN66a6sr5sxVO19uRua34tw+K0SekG7UZwW8QWxiPHF5zxIhzepHUmwTzJAnM9Bw3jgpKZdCx
7mi4DNcT/rCgMrvYD/D6iQJO3g4b3gjoF29E5rbSNQKviDNMGwA4oDdJzZOGDSBXzQAVQFcpKton
NSCzleoCKlQ1Q7qTi6YyOAl+m1+eBuGAMABg5eHLZyPIn3K9rki9+Pnja3atyLjEwWOdZI33HS+X
RA3ErPG+Jaslz1Bqn5SqaxCmpQwBSbLIjRxVp46oXCkXgJaGB3Mzi8UlpmXkMrrRQJAu+PmjHza3
VPtuHbOsQzPndq5nzDorwfNCGid9FP5GLWSvZXey7K90g/cqPZMGHdg41DS5wuuXb3o0qd6TSb7t
jNSll7DW+4CQmU9TtDBLOVduvn5VU/KnFYGJuexAMSY/yQqyNfF0+D26HE26Ysca3oSh6EVhYt3n
lZA7EDsFbPyCLOIacEkiJx1ukYIo2H3/s8WZoYBhU5hlXCtSBMXAt+sYWXkzFFetCgP7fdcR+KMJ
N34upJ+qd/UllhjgTICVEC9YTqCf7ovCfC1JE0Y7n/koVSZ46PcDYbPoFVd3/ehixycOjWhXQBx+
/jHyv+tW4r60iUvc/gnSv3CA1qz6mU1b7oaV4g+2/6j0ungP8PQwQKPx+yfqSQcKHveazos4yJMT
wKV8qgmHyPjxyS98LPIi69X+Q8mbSl3wuU/odswiaC3Huj6nJmT/BFYwF6Lay5uFKcNp7EnSNxPz
MnCOEUvtA8dt0XhFtuwm97Bh7Z7iIT7P7lCsRSY7dm2h9OTjlfAK60G+31vdwH+TPyVn1UFKQGTk
v/qzVPAmyzXXYabrDGMg+eHD6GWleJj1ToJdblPVh1WLN/VOvXmRrDEgp27rFQtg2hfVPhnEmNdo
wXNjUeY4intO5RlN0Y/zHFlgeGGWtvMd48oV/SI40WONmU0Q2p6DvCrEwEqVxK65Gfax53Ag19t8
vlzLvUOv/omHz4SfXrnhTA4wz30tBdua/OsPT1yotQvZLiWtX0ToHuWVeWc8Qfk6ZWMgQxqKq9P0
k3vuqdjSp5Mvgdu1EYhxJ8biIrTsqcp4amWhi+LGhsU5GJ/4SeXJ5E/95Lup84IMyCSY4eQr3bOj
V39+raUyRsq3jKkjF4iWDZO6igjNTzAcKn0jow69EMzgmCOPEUJ/ZM+J/NndEGtJY2ktF5FU/mlv
FSf2D19wEsa/vp7zIpDpCCWnAhnwZNt2dxEmAx4U7NYz5jToVYSV5akMu+WrQxS7BGCeqgajyT60
eljrOomx2oMi+DJOBZj3nEcBR2oznWOyWd0oUK4HpYj583umvQm6zRtHMkkaKFxshMPoP3aNAAs0
oTPYgQTYCg1G5+iPlEg76ScoEoAwMmxU6yUCqrfvQWcW9fIpH3dYwok59qv/upNt9nai8Zucx/Fz
e4SjB/3lO8FStaCkaQpoT2bU9M3tnATMGSPvgQUTRi8vQdCopgpK5ajJoXr3tkqpOROfKzuUJjCl
CNZy/xhOx0IF8kqXUy+tkYlYrb37z8HzdlBbXjZJdlsgYv0yYcPdgqKHvqI95ZpC1SGO0cTlYEKZ
4/grJg3WEJy5JD7slpkpcFK+Gv+tJEvdFzVYm0pj61KYqR4ougmKAXL7RnsZPCHgnMF8sJ5ws5Sn
BhqDXsYNRZlyKopRE5YObioCAfqZweu9e57lzQzYctZE+5vlon9oHr9TFr/qKUKv/pbs8HCMkmfS
pBdS0NpppnR2Zb1nkJS2euQ3S//xeIlHsry2JqXDObAmyVwsE1fZj5/LK/jNTV6NDnWeVzsI9cpx
mmOmSlG6W2SmIYpi1IFPyfxQIqe0OMiDHvDDhIj0VS4Vz5ZbVzJh1ICL6jGOK+wn6vY0hVMjf2SY
JC4FXlrR5EISsbFTdcjXxYPsZvROijjY/irbL3CCArAVpeTfbYKX/mc/+Kw5Q3bVIsAhkzucCXi4
TrEhn550yboQwjAPWliyO5prweQ5yeKId5WUMCFNJUJOtfoPKo7o8SOrKazbGnLEm9+VLkSHa/OA
uF5YHs3fd33m9vzpDhS63LsYVVmrzQNRMY8Wx1iIgrRdvsPOFS53W+p7wodHtOe4vdVAx9APx28t
WNJh7Mh0oU8wFiNyOkdddyWtFmfZiqqt3SDQ62WnpDVFprnbGEHVDkHIN9L4f4gLxcnC6geJy3TH
r8zWguWeB2Iaf8jZY8/nlR+fRSGnCufff3bWjqLYIK/v5WLm3A4RMG/+6Vump5isJtuisED6DzDV
E+JkIW9wgw6BASXxrx3FInQNnSged05uh2KgiA6VVrw8DYO/8slcRPVfjRxXuOe9ReJvzkeggASp
ocJUJJt3fN7FRMgCIvOYpPT/uE/TAu1OHrf/uuRX5JIGJdjoIwydS+iJvN122O6jB/6MU5rW3kgD
uPvlohLNDRqPTFDi87ADEWYkwOE60mXpqKgBkgRzEmqxdrej+Ke/WfG0/AFjBs2X5LJ1s6bOLHc1
mjGC5OZ2WNO2Xgru8kxWR84DiFwEISh4JHvk0tgc2AmxbndET6Tqr0c3DQ8WfjbbvRQIv/fl6R0x
qA/UQyGMmKuyt4dCJfEog/iAEaFA74FNo0nN/dDFq0/w2wr2zwigjdF64QiMHlIfaHAd1rCHiu/6
mG9f/KUi9b3prR5DriJXzevXAmWRFTk+GBt/PDPHl0T0AbX0CsaO27YMNsl1T5O+I0Nq9kHwXmER
y9fPEt5eE9d050h4VvnDgh2cTrtWkNu5kNmpbjKgCKZMhR2dhIc4Y03roUZPNcLJPS9T+iaxRCsa
F0FbXIiW4kdMJw0yCgVJp7VFYTnGYyORbbUqQRwZDVFKvkRGGZ6kSij3mT3L5S2SGlyO/KNwjwUt
kMKID19zGZR1TVMuTrxWLpJTT4FKhEdejvHZIcjoD/p0rVbPQWGWppcxuDtdzdop0SIQ2UsFw987
vLDFwuupyrsKu4fKDn9yywHQrP3+qSaZuv+ikRZJkjFuLR9XxYduDnDZY4DAIREWQ2x3YSchapk3
jxI8442HpKJVkt5yCop5h9WLzIOrJc+9C0VLZ1svGVqjZcNLMsEVJq7zn2WusvdnzwhZIqoUJW/A
Ol3fr5WwjAEGTu9WMjL62gZzMESAg6W9NIimsc03PVCLo2SwnLTXzJiIgrpH1PAv8kDTuOo96W8P
2KSF8sZ/N4KvQG1ocRdvZDLfyJJqXBJOTbt3NdoADPG+LcP+vobnxrgRQLjXfHKygJlWDiAdwEEV
ZWQD5BZe2srUntfEXkG1lIUP9BZCqYnIY5pjYz9sJDC6gPwxIzqRRo5OTyyUHugkC2qeJOGoiV3B
nhRm60QjzEoeYNlFcJKUREJnbuI3WSxDyAiAtm+gF/uSzhYKMzms6p1nbzhQUE4hniScvW9tfOAJ
UAallDC6nd5l66xoXBnN8TzMm4z482rwVLgNGjEgcLX627+g2mXG6gGzZc4WbEQ0phCTM0QetqY6
XhH5bDU5YN3gSnn+zSsET+fdgQy2LC6Nh+mtckwwtWn2HGVJLxtcGmTLdehQWkcD3sCPHlqIe4oK
NCeDqX5swPpjsupwPxYiVx43LLYw76P+eRC6LJg3SKi6w/fPNNm8khkx7UJ8qcEeU/UcYoo53yX2
z1Pgqu8arEgzDsUYMzl+UkRVgppvV8alBnYB/9IvZl15NIwYDp1jlQg3an1ulij9Gly3+lUhKYLb
sOxmpvAeS5zTDDlBTYqcRj9H+Ribl5w3CVl4/yo56clKiv8HCcNCOhWefkgtiAMHum/jH/pp/q5J
4+zWrWErrnVEjJnOo9gn/l5SuNt6RO2eYALa01xBy+ijyCV2d4W2pEATilx6dPgP563AxF8GX/kt
NtbqgfvtVSt5akaOOy+g8dBAhPBPv7lWEY+VZQBcx40VNUjTgBfcsPvsmfsEYEpdJ27+7N/jCk+Q
5BnXYiVxPWEYNSu592cFvs5/eV71EEpeAG1ZXDtg2wLIt8TD1dvCp9dRhZ5cdIRS27OjDBvUMq85
Of0A6QfD2l+qhC05qv6PPzWrJ8YiX0MLOvk+nXfo8Ndf4XLcBa6zcrP9hdW/2I9tips8sylM/NS2
cSrItZJ5CeZNCcTHvqfcf9n6y5ftwaJztGsTMLCafn4XaAtHymwdvJL9vj1NNXLZ4i4OzO2MuJTJ
+N1fVAXBMQOEIVTHOkfZ7a8mIgotQ3IBQuBQexPys/Va5JepWMpz2NweuC0q8k9pY13J6kzUtx/9
JcZ598xVzpUIcb8XtrRAfMdUn3OXPPFN+TPerYHwOdEXBLaGYIeLbbTS/2xhPKA9fqDOrRXMDEC3
OYyLpT5npKGdujFwWO4/3nxGTLkaY91KHEQinGOabesxrpei/xFmDHW06/4pN++w0H+obkVPvpat
36Qq8Ib6Rsd9RWCrv+nFjgmpIYhPwt5mE/VOK+4vytVvnhWK7lDIM6HmEet2As6ugZf9qbqR1meJ
c6RKQ6u+A9PkCSMKF2lo1DKn81Hk3ZCa3v3H0mHnSZCYMM5jRzpXhdChGdkAM2PrdOslxcIhJM8U
6fq3vv2Cy7wMm9spgo2AYcNDspA7Iq+eyKLLLcFSneoo3zB1lEs4PyJVl7eTr1xBuMRnA2Z4RvuL
Tn525iVtohWZtK7nvGmT5i7EONiYj4fD3BRsfVl5eugfSg9KKt9iP1ogdprmpk7iL5YgPlpFhznP
IKOSH2cvwjzqRCAsyK+rI2jpRVdfoGNy2BhZq1ZbQpDXPni1NrtSPflp273WGJ5kEBAKNjrZxrG2
gddhxAy2MTJzwc13hPwZALCLLgrxbOdtMfjsaplNbUlQ6P3RJtDyB3/BgPNVGgPF7hlN1Mt1KnB9
REH7K5tvbJIw0KWfX1a79Z9WSrs4FAH5s++cfSmUUWT09FHZWpo9xI89qNqp6VBcsoSiWl7eQPfr
Xih/1nvgU6p2oYj5vQKOOujaXuS9PU120p0zFhV74CGLTCPOW04Mr6xIhaSDMAIehdTcOzcakQBq
flcsX+nhUtnVZG7eeq/HrBt53W70nSlXsh4HEEm+YjPJVBzAO+5mCu1ZW4ZFmX8XAQGk5TmPG5Vm
xGLfwrV2j2ep1yk0RduEKdHzoYM0kb5ujoyLZkkIqsm57MDCEtCJDMJMp7v9Td0tXVxFhNEuwZFj
r17wBxWBVHKFBoa6OxqqWr5PtMcjk/0T2Zou57r4bN+IXh6+PXiysl7x90VYyu39Z4qFjgp5Wsji
ZkRvBnqX4TOmmukoX35WmQLR60mHgW/LGHLpCbEI55AyxrdCgfkcs32xjshMSNhmZR4FQTtOIVWd
Hr1/TepVAz1JBlU997H/QtC/LZ6PWlhsoWPh2lmleQR9YyxFRIQADRvDk7EkaSK6GJBpnPVMQzxT
/Mmzo8Y+mYFEWci6Nc1PkYvUsQHzQGUboe7nrJDL5lyFokcnEXSo5jG7GzrW9R6nXC5PHP2yxrc1
JNZ0O5iQMt0grTxcp2lxI2JeyCfO9m5/ep+gW+tFNxG1a2crLqxT2rdah5p/NaqVs2Ny5PF0/nOe
6nlTlbd94DyiCLnBBVHXnAM7pdazMLtaaBDkDFYkgZTUnOSp2v0vgB111dc50yP7hws57jz7ZNGC
89mQylW8nZnGwNKJTkuWxjvf33iOJwCs95k6ILOi4pHM2Vp7oOr+y6++JZStySeuilFtiony4tdv
A+QCNCFa71mNPlKXkfU+x0NW6RWQs7gkDwHQsGSwBQJ+xyOmE7OQ9kDs97CC99qEA8/W4rAyOfwE
1iuKZxFPZPCoMo9TUni9mjgINj8NhTekk8j7S5MZLFoYtXL20ABQZOymIwc16A4on56TXy3outlc
Q96OgkGdbIcMVkxGJQAmff36XRAcZadRecniK/x8AsG7JDAKZRb9MX+MU54Z52RqeT5S3olcdoNp
bpwFfbL2azpBsWlQW5dFxymkuVSpU5dBsQon9Lmu4ajByWYDMi3Uz5qQ1LaC93Y1xK+dV5qKpe5u
SLNMh9p3sSqbWHuDxa5a+49NCMK5ERLC8nReBQbwz6T9+v3lSyy0+KsaLFw5G8wIZ+tAAQtZEDII
nHGkkGpRXr09K20272pl1oWyANdMzb/PeDuHwAh2RqHjgNREk+CSFEXlWQqhRfsxm9ygFt4CgYSy
tvx0vGj6/2rGhflSww3JYXD2M+E5iFCL5iDVgHkd/s6f8mEJdk2VciaJEiwb6E5DwNQLVoMYyPy1
hPYLjtc06kpe1jZ51zqR9lTb8HdN5EMDRRKFeachxFTEwC1bYrdFmDn9yw9LKIOqWzCc7ELrQ/21
u/fRB0a+LEdi5zDP00qR1uyUioegmptP0iHZU1/F/kI8PGWr3c/soFmR6wlejToYpf0cb3Jvg5n1
LCBFrcfoX+JqnOA9+7SD3bAHMv0Ueh46armwc4shvwgAfqiM8gMjZDDRvDDMCCRVrIj5DNQGWyfS
xN7jKvAYoFuPfZK6oMLtnhdmaqraMaRnibDfeWF0P9gyI8Cumv1Qe4rgWKIUywyK4O7sFj5nrJRX
7U80xK8XsdRgIQr9HZ5o2fgaFCTC+AGkb/1cunGmI3DJrT52TD37AQGLuG1EuiO3/R+4OLJlp1EA
I5bF/r/C7cmRHqhCvcSItQTodj4boDoVvtxUjt3dL3/lwst5Qy/XRF923bscDMo8TxgreZkQPJKk
PcwJhG3z17MwSDUSof7aQaN8POK5maokX03xugqZCR/uAqQGl/NGsBmF+L6xu6G+T5JYy/CfbZzW
ANudgzDer8zMmwDitJIFSLktiRqJ/T2XTbo3WTFSl25gV8FiUFr3l5pIGrwmyiR/XRCHH/u7QtoM
7p27r5boMVnRGaMA0gX6QIv43MzYQiFfeGp8g/AbU/nRgnh5kr4F4OGMPXgmINo9GAZHWb85vtcd
9cVSO1r/GCcbMZq0l5BHkE80+wOfFQTUOTVIPWcXcKGpvE13vIua5+zEXq+k0ZjUw0k/tGvtZXS6
xq6+tl/svoRXNc/iMwO8Nx7wmpuBsmoAg7xGcDuaW7ewmuLZhVYQAyl42YLb/dlR24/ZFh6yhQbF
O0eHVmOdtPj94n3jdAIztu40Lz/r58kdn3SorKtGQ+ZYHgo/SP0UlshyhpF0tQxm1LCuWBREQt/u
HZmyon1Mei8wxT3aY3Q0v4Hn62LEnmgEboowE+K1NFZkDQ8/OrmposEoSreYMZJQsPPjWO9/B5uJ
8y4cA33yYy6xF6eSowjlmh4dSKvfT9u8uXkcQxkaohAVarAVncuXiVQfn6Awr+8HR47lz/vKubOY
2Sti6w7gZu/U2n0EEpKcxAppbRCj1UBPDiV5RS5aaceqP+ThAES7ITum2LYYG/PQy5Z/neHKGkQ9
tGD/bBNF6yVJX+jhqvDf1lAiLRJeAcOZzTRAVshF43fruKvTF51fLVbEVPVFODd9s4l4mEyF7pzj
CFRluWZiiwHIMaFOx21na7A52LCHuiJg3fzak+JP0+O+4g8V3Vj0v3cCvwjPBZ0rwVrKJd3SjOqb
Rhge1BejKTakGJ7IBWH5Yb0FKn5o496j1dSNKhOSj8lV+YdBxfIstlxUfVnxoS0tLsuhA+jDQu83
LrkuOQVGh54bQ9gTO4IaKGB45W+OaZfHGVOQmDJE6i/wHFjAjAL9Yo5jUtkRGMJ4hxdMcR16YEcp
7xEyMcNyOOJ/zUP9OyFj/Vo0o6UzsBojLV3WT8Ru9WmjYPPyhzkLjTik5mncC6cVxZOoJjrTWXUJ
C3NX8AnCa01eznQxw1gHoI8Y4DRaYt5TEx1Ke01YTPiPkHfVvRR6ehVDqhG5vUjeEJ8b9VfrkOMc
4gQ9swkPLRUdtSU6ZXpq2peZzGk0wuiftygdJRJG91SdccdV0jV/p5WjeozMPrM8oLshTGfb/L3Y
vzkk34a1wyU3IVTI3e1CTX2LrQfU5bR3btn4rs9ENMArs6ENJaMHJufOyQO1/1yO+1uRKQOZH2kI
6jSpECot+3REKJXlJpV+LgEqPQmtJIU7yAHzXEO0ID3uuHbdhwY5mY8vXUgVI+NmU/FQlM5UAm84
YSeT52WNJ4lST8DGnQfzkc8CONmXM1gavC2k6pjBF9xS6v7TIGqUo7VwQfOL5bN0cIJooSkcFC6e
CKp4SqKOhpBNATvBfbEWc+zJYm8Y5l+dypK/ltealrSm/qGw7ZQ1UUnjiUhDyxG/G5w/7TgFMcnC
QAN0+25i9Ny92GBYNZrnlSGAalhY90AjVlGYOepAUCRrLlPj907n4HBVVPchgRgD4INbT76r07cu
LzumacGa6msO+jBwm6A14iD2sa0RUvwF5Su/WI2jCcP2GkhA8NfEq0LOwe/ZyJAoLQuuEs9cxfGp
sIgfhqQc/zzGoXFrZUl46r6ExMqjibyPTy3d1XqA2ZosEfvFgUOdjZBc3wZjGIpNAc9f1vMLKXCC
+LPDnHOaJJCqJG0+xeWHEGkDIAVMNtMhg1Y9JuvoxzBA4XIw/cVToJPPBG/wSHWR2JHdoL+yHkNL
rlH8oFtEg4Yj3XlO47Tl6gFvA00Sxslm3WxPB9qdOmW9NLmiR7jVe4dbuHEMtt4uhRT36j72tLS5
M2dAuJ+Sdk3BDRQLKctJXIdzP4Ln7EwCyW7R9Nl2+E8mdUf2jqFHhbC3XFJE5ZIrziDwyexSzK3V
x2U3/SpDuzGTbOcrKtBzrn1vwn82TzOnZSYgPpKnya5BhX1x5gdH/3FopLgDm5nXj6u3GCeWQWsm
Ypwx21oDscBVVBKz3LEx7ybRsFIeoxutABX1vHJtGQNdDMvZ/S6rSZn+7bKvDQb5C6izKTyIdiLJ
w3uslnH1AK8ol7OV+LJejLvsOjFJL9/F52RmXOGJPiIiXwD9G/xgpmSjcxktzCQIz5mRENs+ud7j
75UT4lci81ep6VcqqQVoQw4Pa2vq96TRfWYoI9YXsjMmAmYNhab2uVn0lXAelLwq5eVuXyBmpmCh
vInnnSV0W9zIjodzTz3k9wZVEhDoo0EzXOnbp4bGSC7Z4FBUp5XiVFCESLBzNBROFsRI52SRkBBD
weqGj3UUYPRw0JEFQcPUG4q1d31MhK/D6b34MRcTUnF9TkzgQRAlOuB3svHwvJwC1u6G+EQLrRjy
cRc8TiA4V5Phy0btJGFVVL1AEcirKrDRSD3jzV5VS71T8Oi02b4BBM4XZ9W6yhtcmABVYYYSw7jj
0JPK0DNK5tOp8EfnXamJeG/Ifd/PAb0MrR+SvLc7N4W7IcTzhdm66twE4c/xtY4H297L4TzBe7uT
28UH0RGlxmerCwxGfqryVlaxcGSlfAD6zm3M0d0JfmNNx3AByNfAocBcS5XhlXPHXe2FZK5caqzG
ENGFUNF0zxmRky6mXmg/ZBMyWbSAuKT8N909uHyMilqhwup7vKBPcj1XSOuhCsbL7Yuf1h5g9bzl
PRFaQzB7Vb1y2tlE+eM9s9jh2aQir+z/wj906C2KosozIY6faa4W6e3BZ1J9IWQzzf4RBwpdmKbb
Biq2JvlEq7HgPIxsl8s+TOFfb9QH40siaMrfO2JnmOwQjvFTtjhwjV8ZcKGfYLvP1HPt07+KkLGl
E5PZA0XAVL6EsBU4scDOYpo3ll9AL5ZRariusiuPTDVnmqJGFw2rvLAx6brE6OYhAHewLxtB0A+I
T9kO6TPWr8Ig8sBMICbwhCG7b9jYZYW/sBIrI93zcXa/xRLZtNMHoXCR0UV/XZISjUd5dh9Bl0tG
L0VRtSQQMfRUlVcIU/2Jp70EmOMsw6UIcwtjsG5sieVDPO/g5kNXtE4kN6MHr5sKBIsqmFv0uJUe
N79O+q2VUpiEJRz0UWIihK9X0XSdJnwDH7MRnA57kFQ3aLqQxVhQmbOWp5sWJtm0qOEuZldt8d/Z
DcEYQWHPLxIcG37bN2BOlFu1CfcHrlnROITDbqnRPM7kCG9+M9GyVy/wYgazXhpJkeggAYmNOI+y
iWB9q32tOiAYiAC7dz5RAUe8z8HTCxya9VBTe6ipdzXeeW0tsFJ40+X8tAshCAf5/Twt1WO/sEuk
Cq+oKU7N9RAvNkGBim0AvyhsATaIjJbCr26KLvXtctZM1FO1XBmwyHvghYNh4nNZGpHtkwoGeU74
HVWtU6hL8IhM1qZJI6dbeKgn/1TClago1DfIzmz4B1u1Ks5sSt34AWtjcRRXraytiW/3KISeRuRZ
OOJWXinRsOXdmOsvqT8x8PXGQYq/QxYGRAK0d9AL6JWNjXgbyvI5yzJsIIPQIpn9GJQV2pjqPj+9
krGJh5luuay1vf936Pi60qOiMCvt3zPqWiFdtnKgbN+x1xG2XN8fhKz/MfmSN4CAeBbAjix8eJrF
MYdea5+4tVRyS4+QzgoE+iRBBU0slBFAVGiS+23uwcXsE+IOrI/2xEdKk6f196SNCIxfg1I/femM
aRDjHuGrbMv1Vt+6eauE50ATMA836uMpv2teZrA7VA0Qx3N2behWg5WLUt5xQMFzbe9vr973sty3
LegnQDIPERRh3OUYjGLG+HFZjmEWbUsLn9/9tw/M2ZntKHjyBAzrfuOCryxt47wr5kpUJHshDT2p
YWgJdYShkq6wiwYWNZHZOjZdXKDV9rUcMXgASkqUAwX3ijCeM6DpO1L0SPgBRHJ2ovBlesUVAcdJ
Q/35ydaCoYTIk/POtA/FaZZde8pwipQ8DcGoRgnxZWCmicJiGJLJgZZ9THVYdPbcRw2ukLKl446U
a8rnruDgE8ExwrnEcAaCzZJr4Q+s5Ico8OclDsK8Gk8winP89Fupi3VdVlZnWxop7Jwt6C3L1/Gq
V5PdV6E1MdQI7yTMjyEyB2sTMyGw7JlEaA4PsymKAFScKm5UDoj/Y5VmNuCA2cNkskJciLO6sk6l
K4MNaGiQP5PCeX9KvEPKKkZ2AUjYSWwjyHHpSSJKVHxVKfpWkbZN6bAG1r0IhOL+/4kOno31lZEJ
z/eqkheU2FQSxtGuRrXLWr9fvnsWJLnmA1oPBgLNVoEhwyR7DZlfkj1Bv28XoBOMMem+TFsaOIxH
d4u2h9eL6QRZKoXFFIZtaB3ra2s1FLhTtF31BG87spcYi4UVKHULWuuBCDyix+fmeDJacmj50VeW
ZbmTT2Qj4DxoPFA6pTriVTKc3H9MdeS9ivCTRaCVVbDPmqKlnWxmp5TDkI5rsXqKvCr7/RAmaEBX
Gg6p7hquUtbt7Av5UtS7UpJQiOZ9Hf4vzKlF2T4IpI/Wi0YLkLSl4B5Sh45kO/3ljotQIb3t9vW/
8fJMXGhQ08jGuQQy9bBAjcwHPN5LmY6P8wZwQFLLhsC3stw0zRI1hR3ri4JLpPjz86sXM6vulxYq
XbB4TCr0g6M70bCHXinVZik6AuCd0pUJa75X9tWwIe6kBkmn0QScXnk7TNXgd2cxp6HIJ4IGbfli
XTUQPZuvNaGKZNK6FgGaJN/3NwnyqO/n4Z7Pe7rFqy0jo1L0aBrzjErl4hi0tloH7+4Ay3K9jTJJ
GpERjCX7agJrb7HI0TVuU/WDEEB9pCK0IgqqGggK+9/wAJo8s+XzocGMO4khDeq3mk1NMlXlSumg
jiRSRDrhXVibae0j2W4O7BgJWzYEaczL/KaXDvr+3Law4OfBJaCW+lp9ESUxbtJ8S1JYuxD2pw+r
yj+PH0QZ+hCjrzdfAWw0hJMSKhelcSRZi1te9bBnexi05yEFTE2nAmwQCW6jFdOMG2dTS+a2UAdh
K08MvSqb0fRMB8MXmOi7FPz6e73B1XK4XyVehXkzrc+VfT5aEz7ESxhhqnulCPG1l0DVqZQW3kTM
fih1XgypxqcRbg87tWfBM2rjm1Ft3VgRbQeZeDvooCmqSf/xJzewwXVOJD6RJePoCyV0poeWymZP
4lhwB1rsVyB0p3F7M97b4zSRefTNipiw0O0WltH8hgfIH2ICvktDngCGmjHDqsFCuS+BFACTDk20
5gVdi0pRCyzfd0QP7DeO96jboBrMEDiOit/TsRdHe8x/48GOfYrqkBeg+SEmxl6bDwZPSnQl+N4i
GAqGvhhjc6bSCiBEpZdzmBPglOah1cFgxapT2DV7K8V8z4qi8Uceyww3bshM+j6qQPDHAxKNK9Bl
pgEr9YCm4tjqod1tu7vEknLXCqDpxs5W82x9K6zJEgZMCvMB+nTlb9ySRZ3/MWuWcy+NOpR5s8T+
oGzL79QCzltLGvMyyb11ihxrnn13oiaKNsIbY6NgJFjs276iOb8ymj63jk7o49SNqH/TIobOdcwu
0/1g68tOHrMw7ZFMF/j+ISndOK0hsNcdb5Xptw9FuIFMho+4AOXabOaTqcJZqztNzA9EvCd6jjSv
qYG5lOfbD7WxTJyeBD4PX+ZbuqXuC1KdHy9ehiqDUDAPP3li7QPq9YNikcETc2rDXSp53lV6Wi5k
ELmL6StQvrA/77WbsjB8skB07exStJLiJXIhK12p6JXJe72wfeX33JXninp1bhVCHjtavcxgsVRv
2itKXDP6UXQhTWDNHwKA1dP01UXCUOZprXmMQnUDXgO5nU1iUoHPIeekG8iin3gdc7LeT4jUAEpK
A6Li9qtB+1Cl4Vr4lBo/j8rk9uaI/rhXq4IY5kYGv7wqOGVblJMsM3fR2LFkciCboa92AhNRH2u7
0vZUMIjTPJOyh51Txqr6AXuK75+4PEqcRxHMEa/pYvXTPFAM63r8HNmSEy9t2iKu2NShkLvuco4t
I+ktgu9Z3NC/gwesvf+qHuno9Eg8xMDXtXDWzerj9vTTdiAdD2sHuyHHm9GbLBxcmQ22iv6EK4ey
mraRKNGKdnr5DQmAsJ8GoHzOooZXpCiPItulYy83VgZVErhMGsI9twidtqO7BtH4gQRd48qhkCnt
cbSDlO1PiVCpmgiUGya941nXGU+aThWinAuLyoPxboFbsafl4f+0Bybn8jdqpgKa8H85Nj9x9Vsp
T18/hNkOXEgBZ6PhTRDom7BiWAHjP6spdTLTFL+Ybw+PRxpiplwDHcuZVI+4gduC6EL/QLP74l10
zatqmMzdQM5N7jgMBmGqlHdFj86r30GgESR6hLRFrKxRBJXw85xLezWltNoLhf2a4YnuL8BfoE8Z
1G8PnZGAmrnVzeJxm6UPKndHp/Xix6Vhq9WtUz5KwN4hkNfXzIr1cNvT0R/ZVVGa/3g7swThyhMm
6kF5rj7LUW7Pw97dRE9fJe9CoP0yO7tHZJF5WDZdwfNnc3YW2V4j+PQytHAAH2V508L06FA6hcGY
XJm1sHkr593ayssZKcVIv4JujDAOujgZJ7uK/T/UaKzZWiOCSML7f0tT6DRNP5v0Mcs/LbVZv+ze
sHwitCvGXPC8wQuD6e09QVsRU0cvaVabUv6+mT2N91w2slYXMS/I2nXIlXqVk26P7h2zmsKwC26S
CgiJyGx8YnIutOtO6HZnJrR17ZrBYolJxLYE2CHWZ7NbFq68u7JlcrnhcpDz79oIk3oq9phYPakn
n4lJXQf/kRY138GPIYpnuJDpy6nhkM1oonhfALELgAusrK6FTv0rGlxM0GvUO9ymOK5zzLhOYiS9
r+cpISnSR5liJciDOhbLRGiUaZc7ps+Xcb2/CJoZaY2AKTgEtnpVaIB0mP1yYfMr1q2A3cCzmS2Y
r/IEOi8paHD/4KiYIGn1IClrPacOL/xWEND838TjI5k2LMEPqfAy0velzmKoTNfPXP3vw9Sz6FKp
ZoDaHqG5E4rzIkAl0KpoTrqgmFtKH5yR3knOsXidk1boEFbFHkRh5Q+E9Gq6olQYF4Pq+DYQ4jWh
dHQkgl9LGtdWRc1JkLLiW2VUhiP0awXFUMWdtASzTMyRNx6oWxJUwsq9W6QNiokEoScHmBE38cod
Ej09MoT6C1KJfEFwBC5ClXrSaHkXWT6MzSkvXuuCkvH1GthqLGVWPUe2lf8gBZoZy5igGA5fbbq4
F3HiWfaS/Om05AEAm/r06pfESQpCXL+k/g7FEJ2b3opa9nM0m39eMmAy6WDFcX2Mgjk++bjeCJk/
KA8ZsLbErevmsUQChA5CJ/pmPrLkzP4Sk11ll1UcnxQaQdldP2/izO9kZW3mhNUcJN/wdb3so9MZ
IYpTg/h7XDZ8xKyOUsgeNS83Inq680Ri8dR+YP9EQ6d/07Drp2GC45AA4KMeA7WKqN9hrsuIXXJz
NAO6eqxFnSWr2D5uB61dy0UgAHarRgwOVH7ONNdA7kqqg95t3hfcAdTf3xrpzZEdaRrmOmOde+5F
uO5gbZOZFFpkVs5PZC9nyyIElz4Kc2KKyFz34lDwfLXfkNO1QCC19FrR4KTAR+x44qnNd8bz0O/m
lNY++DOWiDcm4E83giOkVX0of/rXioiu3dgXUciJawTIDJArY1SGagiUQ3R2ljRCGkOc3zcLLUct
GZIk93e0TS5nK0UgfqRwoPWu54DY1CODTrIzleKMB36d0PJCMtO5+bNrR2Nvnw5uvlSy3IIiCsU8
QnCK62Nznp75BjDjDvfw8ZPjC3/bl7qu0opueK8Ykni5OJbAgZ213gbkfnhdIhDmX8bOVM73ip+9
1mtohyITjWCrqMXStekFwMrh92KmRvTfY6xshs0Pt96TCOnEIQSG4wRKSWQiReRAFfm4uG2oGeIn
z3O9DTnSwv6ezFNBS1KsT+qlzp38N1iuV41lzj3puzS0fodZQq8b1/gU4Df9ESlRsYb6KieAc/nw
PS0IP+E2EHCgRys3CIiOrmZhNlU+5OhDmBJ7o9SZXmtJvM0oNf6nM19JYv9uDC8bXm+EPfilzSba
Qq/kZ/R62oGJFRtW1Cy9torSsw2R9dMzvlqehA9cJgGb4MDc1F2li6NdHZH2H6O/CSc5tWv8MqB/
0PmX7PY1EEpABFNjJdAa+U7N7V083F9cIg5gaSficAXr3lmayQzHcPOJ0v+hB/RYVd/knFY21VKd
dxSIz8XajKCbnEoBWcGfJsrHlikK/cjSjqChARb09Q1gAR7rtvwiRC0TIcwsevD7cTaM050em9/x
kxAzgyZF+s5LcciFAqSz50YsH+Bur22FElqsWtN5l9hjsbj9gdFJPZPl1cTQWX47G3BJqZh1GMOf
X3H5x2C2UBNaAuSILqCVOY53gxd+GL36XwFefGPhsiNUApD0R2567uPl4CIiCP0by4LX80v1sBIR
DgimyWaGTv+18CNhcuPHK4MOv1o4Hu2s/qzbRKDnaLWCm4sSGIYpeVZ6x5sza2iw7aIwz5A30ifN
npMGWLOQiM2IKmU+aPXmqUhryijn/fAthDdzkvnjUVoN/sLROdRdsM6UnBs5AgWAVNcHh5AZVd2w
RyCkcBmHW9B5ajhdze1Fs81w8G9aWO4bAfj0X5mwMN8NGtxhVHiSKAkpY7BNEmff3/K5NCq5sMiJ
v2x9CmSSBDuZnNvVJn3NFRIC+Pw/G/jtetbNmYUyVJFLMNiu99X0l09wCIQBdAE9GQXe8zLJ/30M
L5+lAgua4/Z8hmHPStG2EsDjp4Xf+yyoHwm/295yuvfJhcLPadoVmQtV/xn9n47j5H/kEFdnrdCR
jmWFhnjOF4MnJ54GdiGqvqMbhKFTawfRE6NV6kfogRDzzwciWORAZssWmgsoQP6mrQWOJukjZ0Dy
EQwLedlmJJTqVgYiYOKJeLIM/EXPP5Gy0Fvc7ZVhCY7mxA8ScOwz74NKWQkS6cFop6sMtG5WvWbF
yEO0HlPQc5A64TaSlLk0ZiWeBmK9AuaFFeg1ROGz4Bx/uRBbNHW6NPpvT3GBsl+QCJO8jsKVjfWz
nnMDNV6P8l1zZyfCHDd2XqHjAuTNp3kF/P7hDtWY/pGoO+NoggN2mKwkFOVJ9SF1BthXsBxPO9z5
UiDguV5oEM0PyUnRnU78fm/02z3GAunNjM66+jFiWnSA3vipgs0HZs2YfA/Bu4z7VskRNFv/PGfV
7g+aR+f1bExTDKTYciaKNr8Ixk0nmX3P9jkNCYIDZBePCTx4WGnaZGKkc0bfvT7UXS8QX1+s/vRL
YWvvMmyIWL2IRSIKhdKEye2QoC4zFaN7FQxgdSUrtH12Psl/va4qMiXNnNBC7AHsGou7oL+MsnEC
19+ejgu8l2SAloEuAvAj9QMSEJBb7o0NbMCzYL2lkFpk9BLkq21187SKIrtuhc3eYv3EA+0V2OqC
zvGCfqX1XKgnElkvYQ1pNipx5PkX7vTqvtsF0pmmVUis9xeNGdvUIjlKcUrhBBtGsutK0kR7iu6R
ike8wROa0cuRvZhrtTs4BtppZcrO4AlISXxL2PUmB6K+fVhHLXFbwlTBcWUS4mHDcLi5FfkWLFBt
jhghbgcyxetGKM8mIOj7IB8cmEYsSVprNax7h+bTlEhSGSjJLEC12s5JdUhBKWscHUva6vBZatV8
hwoafYV0RgGx8d9wp7cR8MHIAcbeAebAFpevX5BC+pkDQx/BxWMeDtDgrxxENYVmtU3/24IVLKjM
GH7tuzxKzZKBnBnArRSISy6Vo1frK41UxSWiUfb6mzpfP1VKiN+3eJBhPU84ogkDBt9xmzy/7Wvw
E+O6rbuCvnETzmTOAkSUCDE0k435mWSmZYPQ8xe2ukwhIqQFot6YJngJgQZwOa9YkhdQ7iKNKpZG
lCtkxIlo7ZVjzqot/sT7OcyLG2J1pCWRZTXyDCDv/OFhwlqfFt7mbEz4iUdU9qJjjlpMOefb9tyB
EiVIb8AG5TDEcMiUq5ZF0b1trr6vhsOah6hyWb14h1eiNU5HSLT4NhF9+RKQCvYr0n2818mNfR32
1Jc5/CLzrF4teJHM10qHoWspyJjafpAFfm1fND537rNawRoEJy59RGeQUwtNilZ8vwkp3bz21FzC
LTjUnLxatKG0/phphcHOKsc+TPlB5lotMGwbBCSVAf6zDhIuSEFlcQRAklSPTgEClgWCsOnBw64N
ZlyJQsLBhxgDFEZmw/Zm3GaykdB/bCfFzinkPyPxJ9NkyANNNeXUF192ocVOYW1iooYFYmmKqn27
cb3U+NoGOq6MJAaHUaaErAdNKMtVktofslNvPBYLO2fEc22kLIJIDVt9tocyf1JYijyiaLVpC59R
mE125T14TRUlSGq34XVckC3nUzS5v8VjJNF+uJr8zbOPKfe6rOtse0Wa9W5/Ai4o+HgK6dw14ONh
ZskdGDfAXLYVOO21snX6sYFKSxDBkQOnTf6zVm5ZsNxQm9riRpFiJq52lagyGUh5AQMDvolJvwUG
9TFEt869xyqjCrea616jJ1n2f/itlSaEIWH2/DJfln3OtjBouMANKt+xnNLYw+dySwLjg2SlGFJf
4Hwnytlgnv3lST1nG84SU7SaPC7htoOF0KLkaf2H9Ps1qg4DvtvspU/hSsHcGlGrb1lA4eWtyVfZ
6yIpMWmDv0DvjPmC3IxwFIYhdPEjK1bEt9R4FAXU4XI7KkyVbK15xIvrH0yB7H5tkuvRYSmXGxPO
phd3cOu8w8BJ1Nwms1aquwXlXFutpxDfm9ZHOWx2ATHa9WrZyMLh674epyZCOZj3sI4m+5eRe9ep
ttt7A+JXxJDy3CDewFGqAI5F73zNHYjI2YOlNmDRIQPmrsiW9qjQbz6tKrzFK0cHBO5q+Ec36RLN
Mw9Be+Ug0cSSGuhZCmnEFX5KxEs7PTTzqJ3xlP5HWCUp5nz7G70Ka9fjkPISEoIX6FPQtNDACFVo
A8uuQrD2kKUHpWSzeTkAPMVyt27FWfftwbOFHpgK/ifSwH1cT8XGcJopqiQ/zx8UdPYOVmZ+99Up
i5jav50N16L2HXJkLkRg76HJEL1/mzQtIw4zzw7+xDrsn6jBg3NDkQI526qLnp4DKfhfTLNwl4Yo
JYyiE0/9wK1QpFQOIMvMXD977xr0TKeGlu6FE17YibCbZyCNp85f09CiCfgSCY990jDur8zOQTPM
HpEJoeLXGxZsn52laFuyS2F5J1/UmzE/8mb0EYkMP2A8hDWKShhqBEdPRaatfgNZbEsETsnPFPI+
pKZpvheOmCFsMNmL/yUU4Iz5MXsxJbpEPbOg1ckDzFBlfUU93emw0DkIY3Bzfb0f8/g21vCpWiJu
3pBnVLPdAY+g+/GpOOo7isJH4N/IxKnUFeJR3tG0MvwHIRbezgEmibfyVHSq2v5Hbg5t7d8OVkEL
8QFw5ufElGG3rwy8/npju2vSs7DJ20BGQ9CczTBTOXNYlDaZ46/53UXVVIevhkyfaKhxt9VKHLGy
eJnaRHz2nhQap6xRQ90BIQ8oVz83sOUGP6JYB+GuJub2Phoa7xge+Vn3DNkLf9jvpza71ZsIDcrv
h7RXAh8szh//ggenvR3lUBGAwH5HBFPNSen4WpCnk559gvalaJvIFDfnn/Sdr7POCWaqMhJguUuI
o7It4INjopFmXNvgK8QT7tB+V7JevSh46ntsdpKQyJJ+xKp7BU/9d4u5nS/4cn7OexlBmS+ydFgW
o+zUwNGW0orOojc8ze/aEYtxse8UAaS7iHqrFyQlF9Oy3guPYOWzCbLnm68t493YB6RDSLs8pCKl
VdKd6OqBwOCNaTkBgxZqHpcz8cebeGWQScacFAhjvYhZf2cbxfqZaM3PyMkbxCd7JlvMmJFUTWxz
V6wtYrd/0ewGF0yJmlfwjo2e8I2FZoSm0+KRU1VKSowdblCarMRd3LBLK4fEIxl0ctb5Wu3C/oAK
9t2SF6YXYtfQthvyeN9UT13WQkGPdfHNRrFPzYKzJ8bmeBIgVe7KJ9S826HObzJnEsg5MoNVbGjj
GUqho0c8505cACp2f4eZEdvc6jPbu5mxIc3uVHX8sqvRHPsfRwLTiGGzGdBQOZZJ2PrwKyG9YbWo
mwyA+n+W7A0u9l0iq3xz2g3rp1YoTMbE138Wjs4IWVPfUsuK31h3z664IwG65Gvs03Apz8SHn7W3
H5YH5OewE7262SAImh+iT09Dv2VAOi5YDHpplwTCMp8MKDM2O8D4FL8X4jnoljmVB3BiqtA4VlwQ
dwGDsEd0sl8n9qGFl7D+J7u6Ajd7rVSi+YmXTA6Wgrre/8eQXkE3XzB8I/zYaMHf6ymtZs7bOFp/
WpfCWDQnXCxagByyJbLh0THzpZ2hUzmlbuN+TB/joSKMmij5l/HtVbQYGV+taaN6i5GfTEHxdLX/
BqYL3pIf3wZSzfW9KTuAp2VBEkNC63fmvCWS/j+945vuAgedTD0wB2QGGEaCQ3VDLgce8FiKtWj7
ZktfmZ4Yvw8XBmZkeXHcjaBCTVK8wh7vEkW4UCp6bW5BBd2DF6SAr5EKnsLfvQVJnS7oxiGBIsEE
SoA9N4D0hydTzkKxbNcLkNtY9dv3uB2XMqcIRxh++tsjQYNAS2P7VzUwb9LaK5r8GmOaMJDXKpo9
GH68r5j4ahZfK5jXtm+vpHPnmRcSj7N4NAt1Xtfnfw0LrNJfDu7Z7bd5iIoVCdHZeZiGguETELe6
3bMBkRPcJXEbvW6EPqIEgeYcAs8iwY0bQjFvc0Zh0/1dBXG98JNuaR+eKC/4tdB/i9Nfv4Mn7+q7
rK2kmga1dhwJDB6cZxjt+xx7AVpeCFzjGmKrv15pEd2slGWlyTPGzBgSdzyD3zE+m8zIBhFYJ6RX
w6ro460on6z7NsjUsO2yEwcGg54eU2zOy3uZwZE8sYAD3sQK77tdGOw5nf95OcPymrspb3ftNd73
drnSmUjokv4WcylmnFuxsJ6jgPUUYuwL982nMEWZGDZkh4vY02Yu0IOSID8LGA5BG58P5slS5wvD
ji79k3pWyO5OuNjFOwPbOg5W4XQJl1xdsFKUGrBBFElPwnlGFIPVyQ2HFPiXpZss5jmtUOuNcVGn
JcfFKMe1tG8FZvM+aAlV/ZjjadWdm+EPwbQKFD5vNWmModbskGwJ9fdm6VOnpY9ilygnbntx8Odn
0J3VAfyhFmklXxKyk+wJChdyOhC8XnKkHfpXZZy3+KytT275xykxBPEBn3Q/54vlqRCoC6yFScZq
JzvRXMGdr9uAklNPD6Tzi1hLhnlMOfkvnTPBkasO+An91bUNshw+fCZlBgiGuobSedFqTNi8Oewe
0o1r2Sth0t/o5h8s2NdtYkmML6y+1wKprCgOnG5VdNXUS/UwQ0JbQnpSdJZKuuIZ+Y+9Pi/IQoGG
nnJql2Mm1JcgSog1cVx596qjuVEETfcgfEk0fCubQmUVC3iuYgu/Rr7w6oueDIyRQcJ1eo/XWdlV
e7kglXlOATmmUd5hri0tnredVO47YA3xpDDXSapSjEYnQIH7nTM6Jk7k6fI0yTqslvrcfNjGNeJS
KDUYeH7eckthXvsnQgiVPv/6jHgk7FfFhVhIdgHL6eLfMqr9cAjt7KZF+GPQNhx/P7aNnqWrS9gC
gLV+GIZHVr6Q023mgdnU42n7LrioJW9xIJfuwr0rBnAg6n6FlFQKloU6kZfmlewdQ2ROwe1s2ftY
UZc88TVbfLJiEGQR3G7Siup4dgGQJD0caWEt7oPafJs+PjRqMoZmMHUPjn4qCNfjhuiERyw3eGCq
9B9c9sFcChhlzZ98W5O49w3VWJBkmtuITxjul9D6Dlfqj/AtL9OqNDu7+mgLxg59j0tkOXU0HLl/
rvxc4ItMN0wAv/BQ+Xt3VtpDIDZ+NZNINvFZI2pmqZL53JnYAV670znJ+QB034hhTiXGEc9Cn86w
bTgmgyQi1GdzALQgpBPwn7Lgih0CR9M7C4NgQDP4jM0rhRkQIvMeS0/1KhdMjJPuSi0hBhMi/PUu
IR1jl1XJYe8c+OgIImDknqv7w1Zt8QJ0bcwI51M6vfDgFlwDxo7wFmlZZ3W5Ulr4xXXfhJnzKEZM
KaK3lmzahFdI+M1P4zIfuN1Ixzw5fhUNxjp4xGE0FEk+ESIjWxEAaUPEnhRKi9oVz4JsZHJTC2Tr
DRIx2zzqVrQERE3vrITJ56Tf8YB6Dkf5ZFQxF7+QezgooFiRnyZnnxUALXFuJ7NT7dJsIwR1jLvm
A42p22OJHab6fGA/pst4RutU+9Nkfw+ulD7ePpA6LTPzCg/8AzEhgj7vheV/WJT5Jx0ffzDkKpHr
ezgow6b9qcxwE7p46Om2/MOxcLdzzQP051aUarAxI+R2pVXx8llqDC2H+Tz9vCLOEIr2/4z4N5GL
LLJdJrOX/ud4h/gpuvWstop2S8KHInApCVk5G8TpJfW8+C3ksUppzo4OVpWslbksgebicvHtw8at
ogy/jMMUL6mIIOeeoIzmi+N1Kb+8NlJLBjKvdY0kBuW8f0P6y6SNdaMrU0sTquh7j2IJ1Sa+IYpT
8hfq5SLBvlKGB62RjrZ9wCkY06zA5YQZwAbN+z3T8X1jQqE9jLI4a/8eWBs1Mt4YHkzeXk1RzARO
CiWz35HcQR3iX2UHouqZwyN0Tu68y70fel/FywZR6roJNlCwrejtYuf6qyPiCXBo+DgUJsdJ/pIp
HiCoBHJ7s3RrB9c3YSgIWk6AKD2xFZQA/ki7tFvnbYUV97y6PTUwep7xuIlfkGOMOYVXWAWS5pp6
l+k4tP/TfrdIjeDcVFPrzPz5VyDWtK3cxE9Cq6fwniTsDtTeb8RvkRZRM7xJeww+2gzPHPTwQMg2
V8kiqk64IaNkWDXp/P9Dg0EbutpmyiLT2XdVnWPOdewoX9daJVYNik0WpWpDSwPJzDCl+bwEfXGR
6Gja56MUwNHMYjTfKw4tWyLzfAerllzEy+pA0zPB6GLEC02mUmnSA+4j89JMjCD4V0Nb4CT2b6+o
KPecz1Y6GDK0pdWmf5t2yk0lv+ZMLW9cQJdqgxvAPnHUeKcWpEie9DPhwUFjv5YOiHN5xugZibEO
rZlU7nkNbMUYqXoQy7ldtxa4P9vlWFUnV9ITi4cnVGqJ1tVTBzgfWgT3L/VnE4RFKnrQ6dreHZ1R
ATAiYBO2tJZ7+RbpMQBfklcvzPOb4lxC+molACkeTSFQF8q8wBS32LIXrMZRMNbesjLpIR7jQF3m
3DeIW4Kpe59rVEuj3BY1ZNnYMI5A0nG1NoW61w9SZXrVHa6KFy9/Lxx2AXwFY1xQQzfagEJNjcEr
BGToVkNi1oggNzwB1GsLqdiwjX0OgTfnR75lk65r+3Dj/R7ZzsSagRTE38oZ3QkHhPxYl+JFlsIk
GQHrZe1piBRU2uGzSdiRm4i86Ivx0TESy35oPS/llWGFktbMpYmzZGbUxy8WeBfVgQ6PdwuZQadG
B+r4y7pJwm3liTs3nbdagp1pjVHPycWoIOlrECdc31j7yZVd6R55gb+6E1JMTr9qn1+QmHAQeBmj
Sa9OplwaFivvJPWp7sd5j/MFeIiYfL1DI5LJAzYtAAzjFU2TwkTL09TtJrra3/2yBuFopea2CTio
+N7Fs4HoUHv4/0m5qiAdULF9eEKggfKI5i0QXFICAyuR+bl/IRcr+tN6xUo1X0Jb7ERU7N3N4rV4
72pFDPXZcPs+MrO+Eva6p8+bqtoYKkorJsGLtuK3+WHmSIDuyq2oy/tf6EzGednVqoRH3+dmqV7o
tlSq0bOEhrl6gPj6RL8E2K+BoZDv+21IU6XSnkp/zXkYsPyv4hlXKu1JN8G3EWNu2GH89T1ADYSp
7YDM5PQOYuXm4kTflMwiWjbDsbY3Xi8WII7tY1LWNP5VhuWVtKxZsV/AxbLCxODQL7iDhMo9IPY0
heNhaairFlg1vw/OiFpKaSvPRs2xu4fTVf+nyz8oa45tXJ+FFvGW6nLOy2iL81MU/sAiG5MVj88i
g7ULjwrq18Etk6nxrqaoEh5GYrkrua0DpZdaMhZUbb8Gvh1m3nKXbLUYLs4dp1nLL2h4/Scrg87R
YkR300T0Dna0gT4tTVbd7NPRicvp0vc5eVhTJCZiz/Lz991YRkaTnTG3tIysJAbU+O7cB2is1BYF
blKtYrERQQrlcKIkOAPSX5fa0sFC0WQ3rht0SmU3w33KaSI9hdetsyMygvcNK1RADLdecZgNqNJ8
PFQJl8bqqQOdPE2LUH3vIY4SkCTYxr0S9pI6fc4Lh/HNQMgam8FcO/5CsZXbWX9UAiPH/gLwCmVq
vmySq5u9+J/+WydDcOIKVVOzby2i1AAQQHGDO1rCVm/8/cEjvVu21RcFMx/6Qw9rdu1BI8SUzj+4
4pyQXUPPAd1itzmN2ElGXzl9ZLELwbQQvlgFQvJJ48gj0bUL3txI7mvf2jl50gz1eZfTYgP8bMXh
nLtMhCoWkL5xdGJGbOdPTalCkgmcOcoMLxRJQP/WfOsOZLtN8ETswBJG0oyyaHdlbxCTsVlrmC9N
7To/NCUWIyzJ9fnoBed/gy+ZXNObI3nqLNHA3op+8wTmHSRIMpYAnYaOVsxg8o8FPEFfCZLBcWuu
H7TqwMw2UzVHn90ea1fFHJzATAmby+cdY8DNdpiIcDPUxZKqkCH5u7jCRUhTNJe4/IqiYIkxo4cb
vLu7D9qEELCy5VrzQQxVuXKE3uQ9MJeQQSbpWTxm2dQ34H+BRo4km819tkH6iWUEmT7m211T6fgk
SSGjo3lwct6SI2Ef/wD04GOCnJEuk4kk8BmdvcRHXx0t6brwVhNXTbSBetzQpm3uE948HqbTQOpO
AJXJ/IfTdZWvSN/Tjmtg9f2UL0u4cdb/w9iSmSJuc0hTtftryVFUmWfjkZoyHRmy4t+kcNZ7zP+6
hhkIAOzl+zxac/J1EkbebV8U+DUKwTgk2Dg25FXdOt6Nmyf3bfnevzB9XdLtyiWrYE6fi6M34NC6
6/SZO4O4++iyJJph7wJV7wwoJQNaL2OjaAmCTvrY4xVNgbdKTaRnVwXGO2RQ13zNgPMMpg3d5hBZ
QVGOJvNMg8Fes/LtzM7q09+55HpjshOIVwUVz3dR/uEhVqJLbpV8bKAoOUIYqurg3/jCKV2EqclE
RtrgKUG/lK1WJ7SJpwNMwTLcLYBr2Izk07rJU+30gnQvU0QThZLYMMUNtnFZLItg3lJW4B2uH5iF
9lt9wTWGfcuq/jPHYleZ5skkutE7pFkwi/lU5cFAU5qNPYsLdcV8EV5f4HyyUQYgdwaohWExdI7B
RXn2nmkPl7AM1vsKRAZA4TAJgAcrjlAV5a/Cjj9qFr3+mFzeXCWgBIioUKc7zjmPddUX9eAp8i5R
z3MeDZ71/TRoBVtW2FaDf6tKHP4t+G5qVrFxb1p13OQ2tBws0lvtqw/D3BNtI3OTxWKqYx7SaUTh
/jIUUR7fkrXoKcozZdAjtXjuZdCbM1+j8moIYKPB1dGiVVD+g/jCA+ELx8wcUUvYqlXSH18k+qQI
UbKnqoNZC5BEYjG0ncY/cQCAbRnegzGmDOOMp3bCqn10NYRwWN1QGlSm8mQURrq26cay3FRlYWa4
Zy093A3AY3Dkh0dtxVgFtXV0q3Uit+Lp9jFFjt14Myb+c0FzCNa6S7w1Jbitppc53WsvK6Yd4AGR
EQaIbCDu+BJcFpcFNwcafrDcZY5aaQK/aMBq7pnX/J7vRlhv+FpzA3JLDFsjJUJ609oZrvp4V3qI
eULTOEC3DkxNFIxgF1fOMou8C17VVDuF3YeFW4yRiWCbynz8jQ7seayTa+OQJZZPyPCSK9r1DAqS
6tlyKo29a/mfzqJfDcm9IqQHfVHHjC6kb0UxKfR/RqGCSJItpFRs0JlnMawgg/iLEelz3m1VPBKJ
TKFK5tiKFICb9oSFogcMVv+Yp+faLydSG1v7xPQ5TXy7AWnkvPZ1J6AXTrHg2v/FJG/waemGgckp
+ZrNRSGqaoJFRpwzLXD+29sYLwqdQHDC3SA5tGG94pLwT94G0zuKehK2MOtNck6cU0FQMwIQOFEx
R6xUjpoL4yfAf2Ywa+uDfdiupprcFkEItIfhCEXE4YdVUHEgHkUiCUb9w8o11Zsf2506pj0MyFHn
tPYIBEWBLgcmDCVEKCEnEyV1Jzi3KY2B3iAwZjunub45HpSA3b/0QM9DUm4rfaXGXR5LC+o9Fp94
7fxGukkxgqacjpqPaFcwVeoy4sViCxH20EjQOFyv3Ev9cDEaFBsTh5UxAJWXJDcpFoQWhxmZ+Oqm
e/nDVdXoIdZzV0Ok3P7/xQgbbRT1dVB3tIUjQxuuJyH+bcjS2WMEJ59/DOhH80KBxH5E2XNjua9J
eucsmVXs2nD58TI3GVcFRJIL1248aiH7QWgHTGl1tDYUPyKJojvevcrU/mOKFwMtshoYxgpdFtOA
V1A2677FVdTBYjNeh0pCjaiKCINp2f5uoi4ne83efjZOqLQ66jjYpDo0JVGz9n66fP3G4xOXW1zN
zG9YTPmS8WXPTpJkPAJcGnD976C/s408UQQXbVuPzDp4Nnf1uEg3ivNF1b69dzWf1sLqr6eGTDry
SfoaxE5ebwoNSgxMit8orqTPMQuyt545KS6dBq+3ygySpPNtlqIRYEfySWoCTT8GSXz3ZWNTJCRe
+0WCm0+QjOsKDxNC7r+esr05Zulj6tsM6Nx2+tibRSb0nBggQ2tl6TxA4S5vGym4A0aiYUway/LF
q5FCrhb3SyBfq+5ZTsrI74G87Dj2OYud0eoQoLV98kjK2DQb3AwwfAYWwt4kGONWci2krdwwS9dO
dk16EQWbW5jbiAnrZVEKtl5dMq1lTBA5Vp1Usg81CWaGX/xK6h9PsvPIxsU7X/AB43EnhWKbFWVL
+ZeTUfYp17fUJ3LSttuN7WJXBMf0++jh7Fpic6ZzEEvtZnhaBT7z0WVX9SdRl5Hm4cySk+sVVrPa
AC0hmmrk3G1oTFqBb0y7md7mY7RMd9cQaQhytGrD/rZwCYY6F5STbFB15MAwpyIGlTUutFz76l+r
P/ZxxGKFAUYKnUF/+1u6l3DE7nPt5MfzC3wdWk5+9Bai388hRZ6e5LFpbyvcMOSgyJ96FhH7Sqzu
4DTnxoNf9nHQic2QU6twfAWl375Zg/Wq9TMwzc1Qa2YIbXxWnlX7JKG327yYxAtRgYNUvjLxFmZW
0j51nsunT6NSSADninEcI+MPmhh6PNmfD1oVxzv+ZlhU/2lYL5zOnsGrulJlLGcRsIfQa5e0hJsp
j/68pe/5bm0p9P2VzJuUX3WZLoq2ydN65/HTFrPzK5ZoneCjpFz0fGIpDQcBX5cb97df8g4qTkHH
4l3UFk6JS0nNF41Lxh7RaUKF5BJEmV88UyBDrASgvFcvrufr/k0RnsEWfAoCf9+4Y3acv8Ldn1CB
FDqhDxJYkJhijce5JvOJ2/IFO3pdOUB/ShYUIes8kVLXfGcMNzkIvDvH4Qvg0fUnfunwearFN9Uf
YMMZK3pHvB65WVMD+OMuVZJWCfEMBRE2VLs/lMCHlJrpXLevWkWK2JADWFShGLfkgm9EoX9QGpO3
gy8726veGRQNoOB6XitXSyrgoscvD2KjLp7AA6mPXio6IvfzVoRxoWePqN8U2eBi0cDqbkx75qcn
fDhsm/8TscTBdvp/3mLAiPbBw/2udw93Xu4q3kYtWvRceU97ujkESckoNzfzyFvAfPKPfMjXZ+74
PYJmanXsW70iRBDtH5hwAnZmXNJurkD9hwF7b9bIqXZIcC5qAdjYmqlIBwCx/9qOoEtPXA4PI6ja
qpe5Gq/Wa6ixyUDs7C/6FvxSf4FFzRPTIE903fcjEZaBmlVN2oEvN4RrXObscEimfVAzAPmSD1Ek
CoQAgaXpzrXEbk0i6pwz13FfeWMcnrkzvCfPkJiRUcGrvBUBld5yIWUbtWvGGbnTpJNROw+RbmVJ
uIsMTzhPAypzaQLOXO0KlRcVh5ByTBiTh3/urRgt+lQpS57mVUJpFbi5ok95PC9LMkomECRJGai9
AJ/p230wKk7DbwEgv+J82dWsZCxqTtlOAp+0M055YvU6pGZmhCex6oW+gTohnJy8Bu3ySs8nT5bE
9G2F384KBBRvzBJ+e+anTutDVeLPZGhkoptSTeW3aHny+5aB64gWrrgb9j5/MCSV9LISKiC7aCtg
1cWSHmXW28VS4RH0YY/ekGDLgta4G6ndv48yRcc0aVJ+KJg7AJSYrxiefPEikSnRQvZJDCzu3X+S
KDbjrmvlzUQVwZVo60cEp2pwfuKil65FSuDjLsO/tstBnYrFrwCzDEyycfZg1ypclzPIT2YKyOZe
3A/aNcGorD59OEDZuDD6GOzH2kxks+vLAojkIRkLSqVOez45pcg6AK/ijb3HzcmsYFLXDrkHu4ZX
QFyQetR14KYfq0b9td0NrzH81s0u07rVEMpNdhywyvjmX35EJ1SHyXI8BpkrK8295zB5El8JmF1m
TlFslXFO9JVU3UUCqnkqVLqxFoN6/KeC3M+kOCMRN9bvK8EVUVtppzow8CXg5nWfRPzK/mG1eMII
FvIuVIpf6eQDyQnQFYI1S2d6VmMho5VuO+HsMnS60VklKYIpfLvq8vWWbE3qZQqdQHptYT+vuhhD
BnrE6UW6Od+64u76vfWMxbOZDVJg2FedRmcpa1pEEtTRQZSMmNxuThCWkcZNZHimkw458BkzCVN9
Wyg8ZUjeveNwIEIZM3Dh2/o+60uVa7tTCJzL0WKwFkk3YhzWVbvlFvlJmDxxTRNrmtputh6UU9v6
YBLitfiXYySNjUs0lvgifzEtHIEGBcsO27vhEyooQh3VuyPIrzT+zWRko0v1SDHb4vqEIDGT5+4I
IIhKn8R0GFccgCWgNCIwMfXQIN3QKRXyFRCftM/sureQ6ksCqCFPX66IhSzx9aS7rh+Ajg1Lu/PI
f221mAk86GUvTMy7oPl9Ay2pw6FyjlG/IcnUfamNkT7T4QNeFO/C8L14pKFrQ2/9E8lCfLpm5tsM
cnxY0uaS40gh8vExbF0orMeGEF0QxLFJ/OrUSxPBreM7+nr12oHHohqJGUsZDYd+hCAlVPZsH2rR
eIZFUAFtzJzhkMBNoJTMuU2fyiQCsEFMIC4AdlUTYola2qXRbc5FyisN8aJqq0Cz556HlQidhlK2
k3ttYoMXuYS17ogiG1uR5WyrVtM2S0b/Wd8T7fvGmjEZ+YXDeyuHoTwt4YKOPxWhpeWg2x49HLsH
zjWG6Ej6K+fDn4QDyKnxmRKMTLQedl8QZk+U4rHPt2NLZcuHcvoaK//1Kg5VPWHKrrVRDyjVERvm
ygfpqbpckx1tsiC+1DEiB7DLz/jZ6BcqbGkGqvXi6/DgCSooQMmw4dPKe2vpLLCsFTxqWgXwH0o3
ISS9VRm/8mE6qd6d8K5yCkwVSmZoaPDVl7a9WHzbhxs1KweTBm4Ah75+WU3/Wh1b1GMirSVq8HbN
+Eb7lB3xpyLTIjahSHeBLUUwrEN8gD7OgT3NQF+4Pm8OvqcqrWFUfn2DqqHuzDSGSS7Sb0EYS7/v
gusHr/hbO11/++LKxoucgZJ/daQSd1s35w+4u8+vsE+ghmYFK7Iwa/xrVuT/OkE9z9TyB9ljkdfy
aDQ0Wh8898Zar1XaPyHu86RxP3cF0OLk3UWbjTSpo5rS12ixCTCGzpD+Eas5w67dts27XH+xVB3o
NhjCSkXNA5+HvXOskzVxjSCbf6lPPdVvpi8kX51lZbJT22lfupL2y6lR2qlhOEVdqw1KjxBpJ4+I
+hxI3G/lo00uOAVAuKV2IDr0382Cz1JsqRD4/dP5klE+36H/NRK8CD0xp1DWK91BW6qJDRL+ZxZB
MExzj7+nqhY/BnNwsMjClYJJ+70hfXUxsH8jQZB85xl11sFvsLToDmBa1u83Bs6Kd/adS4LEqlZz
aqqA8S/+Ahuk8XFJvZ6S2hTuj29p26lgNFRvhUpLIXSgpcOk4x6sb3e3moH4qZfTSXPBeQPcbQfQ
pRRe3bZ1dfRf8ij37j67R+ZPOPsKB7mzGqI8BGOgvmvtonedd23ghurLdtmQC2z9UpYHCT+XZ1S3
gd1F8tO3WGIuZTHPAMDl7kOGdNxwNqMuPNlB75yVN/ixpqzfvg0BqPWYmR98t9+oiGj0fCS5UcPG
W8pasQWGkngWodea5vm05iGMgnQHXN/RB837ggNiup73ebb5Scqb3Xayq5J25NGvCQvadL9C3191
1dkRAMzqC7nLS121RAXACRCU9xOSace5JnQiETsyrwSHUgTCGU943lzxqfRPm59kSfZdpdBrcLL4
uk6F2xJ6GAUkN7EQb8pj23yG8BA/EZqXuU/YOtJcgvpY9FaVWlGKaq/uIfPaKoPqIbDZTASp0i/M
v3DkCwAtFadSawvyK9dINskSN3j488QGFZ9Kh923GkT/wJNOLKfjUBv7ooEaIqUl66jsDsBzoWYg
lydRgZs48mERcHXfTMd7iUmqQRqHNPTQjC4O+2I+nO5vuYmjZ7+EX8UX2qW/uPhh+y3IERd69RVE
COKhj7RswTw0eoOFnb7CKb1T9jIO4WeIAFScaczWly2+awqqhbvtYSynVcHbEEjwmPRDo29C7zqC
CviFyYVaCxYqCnU2d6k5k2Yw2/DeNmtDB/JSPSp/hbmzXbz931sCxngTVr+enEZp+Gzv5ckdUNub
gngcnlDK01LjqjNcBa1QggC+zNaJChfb8xlAtZ8Fajwa+hsHznmwMURJ6IjDVv98iY5HtVBiWa6F
nvPm5bIMKMKaXe4GZF0n0Q2ySh/BwN3YTETdjZGnSawC3gbEpQviqzLSzpTF4TNEXm9gRK0nShDj
TEBBfNEmyGefia7CXJD3vVHXrY8x83zGWDiXneDG3P6rcWhCahOxcxrbOeeKD6Nt3FLhIc1i1myC
U4Nn38GVnbkilUXMQ3uybzzn470FvzTSXwLkyKi1VHha3Rl4+j6YCEkDzn9geFW1XDuUT4acmiw7
lV18/V+O+JQkBl4kRBjCZ/sVU+Rmgmj+KghSsrkuWh0zIQCtiD0sYxcoLRMb46nTIOimgf8/VkxG
IOf4GX0TTArcHPTlQsJE7FitmQB7PQjkol6/K9HYmiSBE35KWTUkY1g7MuQjhF7UK2EjEYUea1dw
ySxnq9YvPP/DycwMAfrAJTe0NuOD7skQR/Ocpq8bZEMvStVh8Ztxr3i6R5P+rtf1NW3YTWaR749H
mJIoyz0bhlLs4W3njEwL2Reh9ulCwShC9I3lzSDuHmnTu1YyPV0CEnhSieXkYkf76HJbNUxnTWgY
EEXjuh/Tl614scJ+Mm+MpLGgTKCVNI8vT/9ZxBPIx1+XqXIiF0+ZqlLhmNmib7+tIF62tgz/zCu7
sIARuPsMwbk8pCgTC9sQGw7Lacut/iEYv+K+KdfoQA+ATUAOmffReOolyXu2YJkmPAaqzT73VEP1
bUtqqd8rCdbeQzl04DRHZNYUct6/hSfEygq6zlCLfNbznfpBvdTX3gXbBA54R3fqs9X4Fp5uRtjh
6FZ0v2RwmVaxLr9+Ux5BLngmoXN96i8u/xRSWEOAyp0EKl+48rim+UeRNjkHt+7PCQ+xmGBkH5NF
WtUdXBK84kZZ5Za1ybVB/yHV0xhsVZVsKIDNCz3p+hcHEyA+xDa66QM9gLc2opmvcfdliZ51+BLp
38pmIs5Sj0fOK22+KWRjs4kZLAojpOsce+JwVr2Mw3j8lqNTK2Ecub8HB7b2uLNeEAr4wQkVft9+
yH2MXiLO9PFTk3Aw/6BizvlPrHa8xjeYCuZNlo8EJZOTHD/g1kvFBXWj6jbUnQm17Q2azn9MiekD
DMmqytCS0Sl7oSj1LIYUi+c1xkopVRnl3X6ramUcvMt6SOriCkL4X/JoiY0xyYrE3UOStCfene8n
1UrCn9xnUBictT5bIahkea55KtqZBTDjCD/JlHNoehVANXykcK7UOosIk7V21Im81ftcFuRusFTZ
spJwo4Cgs9/u+Qb5drIOiUIB6C/5JXqn9eC9Lg0Up0DWtyXRmQRUZiepRBopvBGUXgB2+7AO3HFl
joN3igpOD4HQwOJlc4Y5IIVJdWyNgHUYlFEQMId6tXlWbTGA60r6E1fEhgKpCc43wXP2JORxiHt+
H6laCXOv5Rus9X/3Cxxc9asWvw+0X73OtSNLzfCSAlov47tnT3t2j2a6jX1CmWnV62HWvArZbyJo
Hx+PjWAA/Aa6jzHBb40SRp7RduDhizaSFE/yWtILAmhpxjBsKgxDkApYPNpk7R4918S+kllvJHyz
kWVPHDoUaUu2zdKgRz7WdUgLJfGEDd7Syk0JoZL3n5Be8dzgvODb+hN/sJ5nLPW5OJ+WsYRFF5f/
C+JVxwXHSuaohFEnpGpltvuEe65DhJQIeNHsnUBb0X27W4mDW+VN9COW5WlqaySBkh2amdGMhr83
oH3lB4NwMy1115emxlL+qGmw36HgYAbVr8XJZHaDFZQOZZu4XSYz/UYL3xU2QfbEVTW7ZotKIsmg
YyvewqA/Gk7FFEvocCLFyECozQs/EJe0iM8yuUQPkgDBJ6HnyBUGqsi1WDOB3j9HF1CLIex9FE6I
Nos52FAd197i8uhPxgCOOUwXT2d8belMsjwHnkfCKxxu9mGvEc934gFIy/N23ThnTG1zGKqyRgVT
kGogQUIO4xnfj1U7g3HmCfwTYICfGuTp4vySZ52PdIxYPTpcEYpk/KQcIQ9O+vk1w8yhP1FqaCop
k2IbJWXatrsK4kSsaEyuUkJv217WYxWKGPLcjqgx6pp3m8TpNHKcflqvTr5cX6wghVzI9Fn6JMY0
tNhdgVs9i5ZoZA8Ytgm1aPM8Mh8VUWcE18Lx6L37koQqHXvs47YXFrQ2jfzCbFXStfSqsBftLcbD
ywrrVSLQq7fhxVxSMoyDFUYaOwqV7B9GA+T05pOs0wXzgs14vTgKhy6RAcmHpan4lvpWT3gPJpWj
CQMhgIGuCNTbbIdkzPYo93Sxub3xD8S3BoNc8bYR0ia9q0O/sKNRpjsGbQRdKlakYgv23lBlUc8P
mAlxW9Bj106l4B+4A+ajF2/zTDvPoG8oG8jNQ5PVWXEyJX3vqkT+h2BZQ5joJqUfGD9zlVnOKja4
2O27ceMlpl3ixYdOQ/rqT7X6hQ1EpuhQSdHG2g4H5nNqHCDKJqqc2J4eAUIUi43479L0wu2tRZhL
kjBDohfdBvxSKYT49zcnV8WglkXO1WG6ZxglAYgIcBXFV/Lir7IPsIuMLHS9nTSd8bvlcULl/uWd
fg3EgZd/TcC0fqVTP7jx37AJxv1wtmIpbCgq2yo4E5AAOLQwyUrli/Qr/ReKGWs1DR9qDXqgPu3U
gIXDZBxzSOQMKRQofdTHvipm/4Z7cOBrxZ4+M7l6lZkmTPC6biSaN9Zex57foxpdheSiQklupYHO
A4rDrZrB+oYj+aW0lFCi7O4L4mUro3Tj0HasUXlXb2mdJotFubxCgal1VrV7oVXWmLObA7orwNeK
YNslsYEcaDE6riXGzCV/G6dRAh0/vNmWgGfdVWdt0xAOcQI1AHCubkl/NrU0dGTXROJi4K4mck90
qbqHPBcvQtyURfmG9kXy4E8buDyh6xYwa3a32ZPE8S+7TqaA2iZlKw1HUkpEqJ/xadp7QP8Ys9uT
9rLRMWbgE9+E6kua1PTz5nFqemTpmslc8Bu2h1KITA5HJlp2hn1ADnM/qJtOyWgM8CYGEswQwe6b
8XKxt9Pmy4mm/e8T01FE5Q6fuXATxb2oLtgf337/gZY5LopgrLL6Fi6gtEle4XReLnB8Yk0ZP+vE
IzuPCC2R4lAmeSfO6MlhMIpXJNkqpE70f6uSg/DaBcw3BkRXQldg0R6pXFthIO4cr6E1obxJSWPd
IP3uKSkvpR/YQ1op/5tKLrUO8zoW7ViR/sPtOFR+6wgjoH3GfoDej+Cd6tAnyOnx3jCMCYFJht11
BCZRbqsGTFprRrKkogtc7IiGnRnqZWcR+w2BJBdB+dRXYriPLxVIuTcvlHBFzk1sDAlW7/SgAS0w
4ZGkdQ2J5QQYxIPq0pCJ/h7R9qeW7sI+iK/UAw7WdCVylAdXSa0Tg74xQ+rE1ZIFnTMIp2TGQs3n
3mFGPHYZo9Kel/pNyixWSoc2P1iW1e0PD63thpWpG+c8szNCPWtjV0aQOIqaYxW8vQgIC75Mw97L
wqEIQJJVH9hSkdKSjUuY0OnVeSCRJ0SpliHAaBI/phyYSVbRU1Yc/ygsKYq3eZQKM04DmQaY4ZK3
YEaalYosiud6P+ndkS7h+f0LjP6javCjwph4dRRmpjM4rQ3AbQL62xp6pLKibhFsae/o7LXNuI8n
wPleuF4mM+oWWmDWEUt9YH7ARqs39OOrtks9ePkuZz+JAs3t1mkggIAPeTnWeg2O5YVkTCt2S2tz
EX22UXPg2M0E8cV8B+VJVudM7bUNkXHnmiy27ntn9yvpNA5P+c+MVPVwHeHCIC9Z8vILsnPMHZpO
RyjimOKutTXZvIbC7phZ8C3F8q45XgiIRits3WlAD/xrRhmdUBLVD7aAhtWi8B/FDINzo8Jgceq/
ZcLYWW6X0gcbCsjpYEc201JnK3uCh9OeDJSjQ1vOIgmt3HZsNOwQ53+biwhJ36bN/si01mUcy9OZ
yd9yJo8VB8mSGVDukwvKsx4OYUz1ajayubAg09e1MImc6K1C+nnxT3nBlmkD8AjaBLgkowfBrr4p
VFonbyC2o32eXNaWmkvTf0Ad4j3U18JluQfrfHCWcOX5FDljYTiaFDz1P4liGWH6hPcTh+14s7zN
WLHM025Ye4nwJl4IV+Ec8QuDJbsEcQbd+I4yU5V7NUmAisLikLdFjiQacDSvI+AJuL8SfDkdYMnY
I+NCApxpo+tcLDG3R+hiwK7rfkVudJ7cmx5OOFLIYlf0tWUhg8soa1SfqK+KdfqmKxY1IgyoYe7h
ue1zHwbh8KiJCFtVol4xz6keLcRB5bGZ4f/uRe6AcwMhQ3UPyjk/zWfaLKKCJeSPwDDahL74pATV
VPpiM8g9r9toHuvO8Kxgb3JrRw78tf9nOj09j2teTCYwcCuTZUG7dlqokdmlJVHEJjj8t8oMK+y3
yyQ8ow4/dU5j++cLKA8TQ5NErtC0hT16W8tIAoJ2zsBLFQJFVCrDUa2HHX+ExM//405eJpW5/gZL
P8caWBjjwwLXP6nIpDXQiLLeM66rrq1hq3jLoK2UvpBiL1BuI73HGmEOY1RmH82Zc2TiV2EPhuY2
ITaLg6WqsN804HlMPqG758hfCG8nriqm7dOHf1kJUcWf+4MYKmh/R9ynN776MSOskdqR7cE41n63
ZssIVJ8Y+XUE7TbJqXHDw/o0RySCqNVawyfjKIyPz5Qbl39ce783ArX8mAK08oMPlLgA0cll6zZJ
LUQKJUmvAjMDY0dacloBMcPjc8elyb7T3c4sr2iHt03lgscSASvV002j/CNILjUuucjFjYn/9n67
4/hukgXPIIetXbeQSAPSSuRy8u6ov64sXr5cXdN3bSSChSlLaHd+3CvV87u+Uw2YuZ4B59P/T/Cg
Ctg0+DOpkT8t+QyrExFFT2jQJ1ZP2OWQgKSnhSB1Ka21R2J+HaRFOSviBA7ylZfiB03H4XSne4+Z
AguWBNUVIzC1Y/PAfiA1Be0T95Gru3phqZyoOmRa7OKRLHcqRC8Q0ntbv6rIoT39G6HNythN7nhw
fsKTxV2/M02o85b1wMQ299RaKAJoKXLCe4p9nmdmcddO8cYNiZOAOH3oRbIUA3mBgmc+P0VJ53JO
5K80X3TOm00CyJtQ6sRDcbVXdEKqgV7NuvkYU+Lmmh/ifqRF9Nf8QahMSmx7lxtumfFKAiAtZ7b0
p+U877zwRv594JEFOhdr6gpPabOUHjKho9YOw9bRf+F5mz768kNoup6bV2As6W+rRoBQ/dezmP86
AfV7GaLi9jID4BaApbK0rFxuqShbEFzNF1dQ/E9zudaGDU3rdIdGs5a6860F1RJzg4EGe71YCZmp
mcrZo5LnuZay6/K/RDyBjSFYeo92TqpmYzlpT0Hgd6VlinNE3EaQ0/+eIKlO2RSEb/1/6CD7d7Xa
aS5i7UuUS/Q3DBGmhR7atx/rJtuBm6AsMVWqHpke9sJoCTOF2SrJ5n767QiYHB4MfU3Ni5q57/jP
1Y5w5VJ+9eIGHU4HrAlLAIiwbiq47bvAA5y2kf1ml0UpJk1JIrwu9sjX5WRrM6BKzL/LNJohLz6O
3SSV1VH3P1JGTQbeXMHmVqOIJkkmp6pIkwDeSuqTfVUCiNP8wOCuxJFmZe1najgJXMDNqPert9Qh
Mt5SJTlPJe634vhMUH7IWFVUHxWBxAuwmOb2PhevPVo/3AtzBppAL0W2Lj3g/m43nxihQmKtMudx
j7cEi6X0zRzb6hvmsRDXmFa847rfrbfZd5mKCcqMC0Pm1sylF/E9U7j4DYBo/hxBl7Ok5TKSJ1uk
KITiSdScYwPggLHufzrlIUPS+9BuhKUMHFrdXIytV0ffCjMige+A3n7HM4b4n5XdTTr/HnWzx0LJ
5LVf2yeqjLJWrZXchfQq4OdO/mti52MuJJHLJYt70woLBrmKRsfQkOXRlFGWT6EkB5NdMNNifaJt
Y786BL9Izic5dZeK0H0biVr/RMIaO05eE7/TvW9rxpXUC6AbsEKb1TOTjCaFtPImy9645l0AZfww
WDdjC/CyVWNA19ZiFn02I0FCjRTpgIFAEorO8/R925JW1U3si1Quzn8gU4eIdmm4jPhk1FNxd9fy
OqX8+wc3Iw6CxORshozAA0irAFAD3O4GWbOPVgBrGnvff5T9+Alv0RygqNXwieDWxJyUuH1rcXuL
//Kpsb0l9Jke0oNILtKTcJ3lD7j1dnNutz8nIFeqjb5uJq3ie85g9eozk3UuaL8hVIWDCF+KrA21
QlJ82OEaBTkfqjNXmp7U6Y+wkNSPykgZe6Hx+NdC8VPL/R8Vv50UN9KDUFBc3xRo8DASDTx8n2sC
/GyoiXR3pAD48fhON5DNwSjjcAKpF5S3ER6rij7YEl6JMTxdszNM+x/1xxideJK3+jV113oOdisd
sz47OXwkwAOoG8We9RmUxEyeEP6WuyghRT32ZSs6pFfj7pUVfk+2gf4TV0qbcGKneRCpqD/v2sK6
JNrHEqi7COTyQ/160KssxO/QNB1/qb30iTMMhzw+0SAIOX7QLBtnxlAxJFL70knKtpCvJGjJbbvR
Ab2mzMVts5NARS+8B9EpEOv87UR+SD6hbHNjbKAEwRgSel442j92/aIMoJVN9AH8OrK6i8eZ0llH
AILo92FIXrX6Dy86mKrtqoHgy1MSNOHGrO8vfbu+8R2KyFAA5kWyL5/RBXEVbMkIIz6SuxxfJ4V4
aaapy7zTT60drvUcT6zRFAQCdSB0tECphPjFqAMXTXlkVyXzQ5U6epLIvZE9zWfl3X1wDYeeKQ3t
9BxQ1j464rfKNEj6ibPgSEbwfTMpyblKrors0vZG2KYz/psFZIGtHeVeCkkkDMN6X80HcQKTnv94
VboxUiI+Wgq7gT0B27X1Mq2foMymBawSTzNdxlxKOD8czxmhZTOfgGydSwZx8g/uPj43P/YFqtHF
36epiWfa3EF/XnKoTYx0J0RzpyGDbxwGWxESAXRjQloLMbgCDkSBifM3s97P+OFh6DVSml+ju7dJ
qbGQ23Yqu8yNtcrenn4fSM1wcNfNyic3Rlrd+rWV1SeHFghQcKcaEYZLYbeB7by+GA0QKMHkUjTM
UDPdPKnkiF482Chancu416st/U3mO9vEGzci2CrzDjTew+vkE2zCQ3r6DZMsU+d7vyjVsGhNJb2B
96ZOeutuZ5TpnQouSase6+Wy5Kk6Jz7wY/r/9e0TUtjoJ2TqGPH4CAAi7gb4gIU3P/iwuTMTUZnj
KLcsbWgGy5PpiJ25eDghiAuN748+n39tt1uRw1UFgADkHXPt0UDhM9yLWtNLylA9OAvyoUKr0zCA
q3ILZIcmlU7y0zSGNyzVnbwzaiNPUz21PdQQwt35Mto8oN0ruotEfkDzQcqkhdEb90qgQH3yIbOh
jNWUwuMJV2jJt0jSBzPyA7gAEDynVCKrshn1DJPyHR5iuTHOo3GM3MsYr9NJuscSb9F5WSDOpFXa
+D5GNYa2mH1JRFPl1SlJjJsDqZ8lU/xrenQpzd5mJ20G/egz8azNQqriimHved3EyD3vZnZcjhSW
dHt7PKEABvupRfvnSz64m43MClJ8fmGWa4JNJae6SRJGFX5zNHUrJkZARaE8WsJSwpUSvH9pZvhU
ECCZGGwi1sq3/dAJWp70Z14mi0X7h/ufwQf5bYgFO6F7ow2qj5Sx76vH+rIKtjLP2G9xJjLMf5+M
ZGleg4UJfb7drfSIUuoATbtuVnN1uFsjSAqe/GfQDBqIPTatYU7mmqc+id2JvEIePxa/0xhNh7J7
O2MaJjdlc3mfYevFzgpomR/DOYxLoxpPdy9sobZbL64G2XsMVHnxDheKo04GtQpI92bc45JLyf0h
q3my4tF1LTaGp6T1EH+TjO0WDjEp/cbJ0QocxlsJBcUmI+gKZKKPB8u6iHhoh9nBFpGwYf1T+Iyj
rMG5SRruQaHoWbMkK5/XAaa2j1TVTPBgC3xCjOH56WJdwN4Se2EajaxdU+9lhLcuneg15ItDeSD1
2G3OViemJjPPzful1hOqvSpHdJBEQztWBNE4FUYIx94pexixqi3gXyG4+p2jiEqJy1bfg1v85DTX
1Vc+rOXcAb05i1Oq2kERV1F1Ee9+d6p5/o3cNEdBtgIs/TvlVo+F62ukH4hfw1+b427khY4qTcjj
hlO5Oh4YGX2mgBWzDjnJoV7y96mvlp4dbi/YzbtGHDsvtoV2LF1WrFzMIzMG8EGP7OvScW3gdL5/
hn6qyNchKkJ5KSUPYU5+GxnNSqxoGeXlcPVYjhlvCa4ypi09qZopk8zsHhcKYDnVMGUlFEojFfKA
GUJnmGktzdh2dSv8mZBYuKMJSpliKyEsdqkrcJ9v79UHsVYpTUYVk6A0EodLABMnA2VYOMfmJKzv
Skw5x+wdCeiPIAMXYzmTvsq2MnNox7gy8uGWsZlbWuQqfquei28bL4VcmD2RJxNtVSgWbE7zJtm/
s7Ny1HIhnThUnp2XdREZwCI47ndyFpjlw0PpUGQp21mH4ado9C0AZJxgHc2upBVIv2UxZnKUNJeA
pD46vbcFXRqyiAC0g8uYb3/SUkD3nTKgI5RTtLG1icnZrSVLi3O6b0zz3eXJeNVxEY6NCGJclkz3
anJqySOGnnME5XldhDMPtrvmAsYvSfEZkP0/5tjFFYB8RvsqV+F3slcueyi0OVfiMBS3gHKitgy8
D3kOEt0fNrVZfZY1pI43AOiwSl5FXQmggBdquqhSz/gHNvyBxSWEPYxOCkejvgvDTCjJXYzTTWtg
Dg8RbzMkoKcA7lrqFxi+00PEVOWw20Xtr2+ZTfDOTjo7FgyD36WS7a04ExSxg81FZNp2bN8pBhiL
UWIzHIRzHuEgy27OBP1DeWjt1lXM2m7XYy2+XTlJ7iOD2Gtz5avtJU7t65S7JVNQFpV5f4PcLdsr
IApfNg+ILSJ/MCmPy+89sm1tLo71YbmMtv9R3hwM6XlepOKDbaBSQkO3NnCHqECO0jZDi4F4VhWq
7msMDyIH0caKsHpHuObtMeT88hhtBQfXqi18R6jHYs/1nFg1XEsPcAkT3UEAgrrSHiVdwqIl3Js6
Oh3qhps4ZJGm6RlkP11gABZNJgwcjqby6qOAj8zkZn60fU8AWZ2inyb8Nc495V/txFM9mlozraNY
YULeOe9ZQO2SHfQ81WKZHUtHJSskiKaQCIhmkbEyahl/BDBur73duAx15LroYrHajLkgQ1FQg34j
gENygXfXWQOhZgYWEIlRSVO0yvkhQtjhTKhaUIYGcuFE2W8+RbfdVRc+zfa0VRySDRX11KBIGgWD
GCcUHXI3AAvkPV8cq72Jq1SdTzCRhnX4vpWvkGoZTsMrmRh+brJ9dzGTYWtfEX+OcYCWoqsw2yrE
NpcjKqKCaWaSsCPdsDEmTDKZ3Ygvo1S778yFBUmyYN7dwIr2mLzSHqjuS/PsQwU1GcM9DXNbWKHd
s9dky6yh3qFYL6O/Txi//R8szPEG/Y57jxs1k1/jEuusSr/7oNJ6QcKHRbh2ZYF5zXLFPWA/hVCf
TKKolyCXq+m4+GL3utxyWMg+fL4LgubSz6mz9n8tKcqVA1xEOtjtuwpWJ6cb5kBY0K4SQKo03E4O
39YkftzIb2KvUDdgpgNS/zaP4YtaNLrjqHGeqkSvH0ICBHTJ+fqOQefkIxHWRYyUHleSVTycw98V
Lf2Pw8Kn1wEDPbNuYQMq99kxQe0HZHqfp9elLzAtZT+MywH7DeBp74rgIPeF31rzLVNZPydONZK1
IRkZzmACiiUo9iKPUfKt3wTVATBcdXgFrfuu0oNetZHJcI0wOU3HQf87yNcAIy2pO9+HTYb5AJIl
3pxKqLB/nSDxJI01G7tLHnbk8qMx9iZNwvKm6XYCAgpi9hj7VILXgvK4zuVvvgT9SZP6QCI5HNu/
IM9X6voOd1UcpIAzUZPyKM6zAMkJiTG+CoPdTFhtZ/6JIyFgaik9FEMB/+WdOdadN6o1k2WTU/rk
coiwuJYmN716n0qAZip17+YAZHmkCuZ2pvQq1xP31wJcqQ4WFbNS+qh5tplh72DICyJ669fgx+77
xCRztS0XsBcNETFSDdliDVfOL81MO7UN2XqlU1HXRVq2FpmyrArFulXkNxpXr2okStygrY++KBBP
ji9LyFUotGl344jy4EWC2dsdX3cqstR8fFMkVgDrB7Vk9nsnTrHzFaj1v9BcU07PaP9snxn1tYNQ
U2pdJkRY7NuU3aX66ZAjgw6PQEtWizMgOD5vvKs8rR1vB2wv4rbDjx91JJnc4lOKeiYPJ6f2OhPE
BzW51Xyarf7GdxkZshgtbHkdcqgzeJtrbmmeE1vGGnpYQZMSSGrFQhQXXKanlrRviBZt3weBo+7U
9WS8Y1BgJbesM11YWplYDRpoeDCHJpu4rO7djO2Qx24zPGYKMl2ltPfXLwB/UJu45zIY4x3kdcFk
D+jHF9AHxIeRrIXNBZp/WTZMZTORr6ZJ+dmmSVZR+6SDo6J+DQiDyGuiLJZBQlNfOR1y18dUmr9f
C3mC6vp9W4Lup6UqXdn/iRjaNVfOrZ/HemmpzyjCJ4d3GYEZ/D48PvQ7+zfXzhBUrs5oAHq63X4a
BRGkUeuDuQ1qv0OYzCG8CKdFkNtajd9+Uv2Gg/nDdhEMPaYzstTlkS95ITNYmAKjPxRaO9+6jQMt
gzupGKhQvn8WTDSsdnxg4pUOsz6w1zDsYBC2T+yEFpDXaAycg2eGBeIo4+5A1BJg2i/inhTmjOLy
p6LaWjhixkn48l8LzLEuVhfD3TQSDg8No6tgFRWwZKuIO29qAurXhCFaJDIBCxanW7z9brdw4NlA
h8bcqcTlYgPAnD87OAdomAtjGF+j9TWHJFbUL4NIqsUTQewqpk3E6lGvPJx4G4catOpG9h2HnhTW
i5qhs+ZlmTpw0WdM2TjQSHUIFDFkItDNflcFav2Rzc3VymjbsHXur630gdYZBBkLdwGU3f5BsT36
7beOtfxeW1jJpo0ieQvxskw9vqXoPhLcO7AL1SlOt8QfqADzTOVUV9Lb0QepmoixZQRpmsJXVKFr
2nirP4BoDX28YqPJW+Cthk6PEOB8vyzKQXSyFaTKNsGEWsHyNEzm3D1lAhJMUGghYSdbXoTzPXOU
teKh+mM1xSy43ievZtMOrfrTPXPZS62JKtlvfqDtdoqMxLzBfG8qAsjN00sIqumyRH3np6LTpquW
WH02HmOGRzE9EzK7npW06gOV+/j1oMwTvdvK4GnYF6Xput0O7YiTyjbpqgLrOezibEZFTPvB5DAj
UacQPMXo22ze0fWzbB8NH8PkP0VpCE1iKPCdOegfy6xR9VKR113Yo68Fev1QvNpOJ+LZut1O+oRk
yJvFak+PPOshNXrVoH6Xob8UgaSo8kMZMdILJtrskP7ODyA2IU/nTZJa/MuOBbdiEleITaXw+zfE
KsmsHpl0FYNtAMbAbU1FMS+mR8GzBbwqZShmNjYxGP2iQKOQZwKZVR1b05LZB+5qZdAYGNIVatya
CtnlnHEfcXNm+n7WKR2TpbFQ8br1EDhR9yW0D6RNqXX4IjS+TEwbTNCvnLRaVOMRyqSOWtVwwI3g
wmqprnZ+lWMEhCtPM/Mz87GvOimfoOyt8XuHpAWugoX/FghdjKePlNEUQmcmkB9x5kqEP1YP9al/
3wFz0upxP31MJzXT4Xjhnr6MzERq7Un2sJyPrNwrn/YiM4dPJDxdoKbyzilmpqkOkNUp7gGge3oE
vW/LyFmqd8aPxl7u0uTv1/3ovSIUlDizkc0/Hkxqmpu2HsfvFiHRGogrL5/HNSg5UNu8V+Uiz0/d
J/PjsEiHEfa25tqidWS7hdVxZ0Id0vmoEoBnnUoZzGEd1rELp+7U1cYmKyJwIHEMhc8PDVyC+FKp
iZ3VAN+U0LWFjmeVZ1AGnU0jhNNc3yxmR61HoMUEAFsHRrGzz2j8fLfsE9qeIMAB/mwhKkqucA41
E5kEBGRCv6QjBagjYUdNvLDIQXv0cVmNRTHrJgUnZC3JAZquXcluYCUTTmUj9QRQQQ1nFkKS628M
uRFd2Xj4IUC+omaLKb8B2O/VgfrldH+LiTykr/j/yUs/A3hUHxA1BvYkwGWcm1WN9ZVx8JY7XJk2
R6j/FqvOtxsPYSr75CAQAyztrCSDtWqSLV/aA9pHrMR6l0wIOxBwx9ejVaz+sOGNSt16mNOUG0r1
gFyHNlwZo1tL0X3GBODOE3M8Hejyf6b9U1erVIV55NJWZ3hnWfM/fscbQm2SlS879o7re0wmIor4
VcSdHNiZXKqEv7LD2Kxj9wmNW4wrkSWyR0Vw/iePjTlPY/NnbwNd1d+FaesV20N/ThISSY5li7x/
0htc24vZ/EUKtr8rNazCbMbyPTVLDn4ezsfMpShlmn2q/nVSBM/NYYimzJv0AH821nEry1IqP7t4
Nr9jDmgO+i7Oxqb+WqquaOFsHKgdFp81p8A2HKwQU9XuRrfkA9Zv9s7ibhv13s4h1kk5yA+vyQ/9
sZjhjMT1rz7vCCSRYi7nUldTYuaeurxYhgFZhb+Layeot2LUiCWV/p9yUy93K610fQ1b00sftwzF
ZXkFB+YZn2SDrm2gexCE7CexhTKY0D+VQWYo9SNoQGF0yT5gIKdMyk4ZYUv3EKaHiiITzPezALgY
cbS6kQ+kXay8sIrmxv2i+nkGfUYnMMgi5MYJ5JDJHK4FlW/hvHF5BCDjL98HxZ/0ccZfTx3FZrAh
FVCCZ2feHD+xdYGlgFi8QXBmkdHQ0WZQOmWtVMmZR3scsUxZZfUE4IAF2FIcJRfB/7MF4/DH3cxH
dCsZlyVqkHaYCvDDmjDuOi04CrpXB5qBJT9KUYF3SH+ndr/jKgk5CPLB2ilPMw2DYl9MrbpNQrd/
jcCboi7fhUHGh4jhqe0jey619vc4qRHMBB9riLYou0ePGHhAK6M02n1krVAUgHDY+ngd145ICORW
Nd5ZMyTZYkLVbowK34khUjCEJJ91IKNik3fB7jZiLgiUMyxURxakYE0ex+StaC4hwjauvDfvsq74
7Eea9MhNp7INiNaHfBJBWetNaRkaPLJQ/FL7sN2XMV6G3OrQklrd5V/Ejqn9afkav5Zc8BiIX/oE
CsasMRA/Jwkh7vTztFpqMfyJvIgioTMVJJA9AVBQC1QJhrex0mBsqAK/zdmaHVERccL0EuzGIryx
xb6QDZ5KZwj+g+/6y6gd4C4+NtSvKRfB1QTFHXjPhs7Lfq82cgbwAfZhJk6nPM73gkymOejckgOz
IJ6mxGuAJ56sYLBAI5jhlIaaQROp6vbwhP/ZwA+EFe2oEN8WILGvSFj7mCibFwItuqiAqLV5q4sl
/zVludY7dN6Jt0+uGG2FY+s/auKc/TWPqZXrr9km7gdMzmX2669maY3RdeA8kbyT0Z8Monj6nHoR
D0f9KxSJ19Zg75VuxNZ4J7lBIR8idobq083DMO3Ot2hAM3w4Fo8TUO52zaHkZeZSTmE8vVhSh+zV
4QS8sln8u8+B9XYC1UxEiAwIIlkLaTSI95T0HlIuLWeGBAQApsIdt504y/owi+yDOYe0D+zDRbfd
JLvUiX7UEtBASavD3hRKlUFw+6CLZbtLTpNMXAfO0aCdOhwMlTs91rjiWUpJc4TFLF+ovBD1v2iF
1SX+g0oR9z6EfCY1g4svgiPAxr9EKqK+Vu1YQkGusgCLDk0IXGg+2xKT501N8RH1Jcbq/dZbJK0Q
EPGK+gs4MbbPX08te1NuVsjig1IIcrVRdTw0m7ezrUvxcMRMmZIQasJeN+QVKRgHUFK4CFl5tdnw
iJse3RIfGz6kACYww9jLQYJaKwLxOQQG3Oe5WaObUYr76d/FacOKKjLyq323nBjHTZkfgzGfXm19
dV6hGNC3aPb35jjcgyg7sRRVhMkxcusFpGRGXaSgw6Qnc8mppNzy4222RQNNgwVsDniU2UR2J9G/
EPDjwWuUWi5I14czlYXZZUiwcFDt8+YD+ilLaxhvlvXBX3rFjIeP53/A0y7ldbTo4F9uXaCOcOq/
KpObCgfYuNSeD9QKLeFH/cj6zbEVIQDMb2JkoLBfiIC2IkA6wjvE+Lp6gLb/JuV4c+WxmleKnfXI
UZ+KW3rnCnGrosH3rjx50E0gN7Mbft563d2sH/UdKJBcpdl8IIWfc2FVQPsXVKmCiV70ZfnfXL8/
j33N3XVE44iDh9tqbdkjawNDL6CI4/RowAScqLaBa5grunmpMZqoWkIzhIO/mQe0w+XfV8VNU1y0
5aORro56eWQL6G5gS1HEdqKzhlZtFYKP9oeAy9tT6flokhFB5LzGTG2VOwMf3P0kYNICMkxOf9Cs
ZdnvVnkBw29/FbZvnIOHo1MmP+qQFtvw90fYv1tAxBXj6y11yo7o+IPSHdJskU3Clreo3aJva9K9
87M7fU9QiuFHCYeHh+/ZC8RARQd3g78CSBRTT2l7bKcriwMAQNuw7dg7tZAK90ww7LkLIs10K26t
+WHiucgjWf++KtUVhKEB4aamvuZC0MdmFIv0adYLsMBrPhR6Zum18LeJTy/2JxeDaRa+rtkEWU39
XZim96rA4mHZz/AJC3X8l3tjXQOS+VsW12vfwPSg/Vm1C4kqEay/E+PH16MVDKT4dONn78Ab1bPz
bggb4RXzSALXFP/j9B3AIpdEllDYolfBr+alciw1tLM0n9Cwr39UHJGQCzrQ1iux1YNdRepLRN25
LcNssbXCH9sLIa7uA7bMtf1Scp1FpiUGpqoSdNxl6Q03dGEUfFu8hso47VR6aN9tuviM6blE1mZV
33CvBS4Baeo22K182YtH+OT+2ntOePxZ7kMnV+OhJuncQ40flqdHJjGM681kcQMYtLOnWyvqDAv6
8/+f/1l28rCs6jvQUR3S3Y5DWhIAgwtL0WwtRMhvx3mbtiu1tU9wWhrS2orRTzr19m5VMhy9fayX
CZfxfw84Xf2TdIvzJkAO6vl3kZ1ls0itEKA9Ipwh+fHgO1FvPA3QZXDo8JD7viARcQZxfdZCnTZs
+SrMs9MBfKUgLNPJu7BpBofQlUgpxH7s4ZWCmbn2AB0r0S+hXJLIraxxuX1hr7kbpUOt7zLbtM+Z
T2wb6pcd+/XGjtlhRNlHhWtYmnPiSRSztfZyIIDmB2oUDSlJaE69fMCwUcMcDLVp89xYsP1o9rAd
yxHS7K+LxOre70xyG9OiL0BGMww66kWDqNA4PLPxr79iYa85/zObHy3tlzF7mOSG7NniZGCovUKW
g6t0gFj4RdfK2fBbwto1hlxJ22maANtIbgdpKo+qhf61l54Tiaf7517BbnVRRg8QzOVh1/LjLvxW
IU1Du5f/vR5zp0myFwiKhoMvQWu8Vwqp/vcCmKQGo33bNHNilXXCEoOyqkzz7Z2p0/KooAdx+wLD
oHKjUoHJUdnGQDz7RdjGGjOXtEydKsruvelTzGjFIsLjhkt1BVn7xngEJNL3qM7MTUmDQCtd9uk1
8uP9vLAWyrXejBgv8/n5BhqkYcG2hFYF9BDLeszWbXBafRgokCb+a09F7qGfhemRc17LOyw3k+LS
aMencSqjOz02wVMq4pZn2o7tznJKdYYC6zRsnhf8hyzoqi+W9SuyftxCLkfF++fQ/k4OdGjRDs70
/zxrjs8pEfu50frp+1yKYnPNohk0PQSlBTEksnKrc/Dqa+Aww1xXgPdFDNNHgKS/PyKNRJI1Bvut
suPtBifOj4pjzVwzQ8iy5ORagweggYhuK4W4L1vA1atIaRT26Xx7prGJeNAKx+PF1YuvoQXOvOhW
cw2Pq7cjEvntrWGg85XbFt3WhR9SnQ1ieILM+oGJSAP6sb1XFNBvMAWIK5F3yhqDzdNnLahwLJdQ
lUGJiTLgyYxjwugs62ohuCr7h6B1zIN68GroA/xFEH2MOxzjbb3fNixPX1uZxboTxfHBCqnY3s9u
I6hkUAjEKvbR2CrkFTMU/euKcXqlz6U1XkUeKcan76QbCXPa9pwHpWNkeV1AMDLLCk9JkNxMYOqx
1nv1/DQ0bQ+LXBr0eH7PH6+bToGaypfGQLDcS19jA9nbHl3L+5U6kBcYED6D7JI6reHhX0gVIlyH
2tCFnXJLGHUCbI6J7csooOoGSFXi8frkMfUL5dzSiJT7MJgRIZMTGdM/t6OLFjHRDITvp6GlTSkS
ndjrBWbA+cCQS5iBqe8CnOUu1w1jcotqybUpKHE8tKiiBW9NYqdwqCk/8SgXKJmNWM34MHUaS4oP
0WEX/EE1nagdQ3qKBxWIn96kffuUSlJxGpGexi3m6MxrFacrzAZFvqaGyRM7qxgU5XSbYUgdQP7k
fcFOLktoInrgxZPwiJS9IhLK23cCh9DBJCKiPnO1cWvRrmW1IcY8uQaR/dN2SJ8YIfO2sy3zKuqI
cnK25/jxhTmm9P9mEQg4nfc3gedLXbRNrHCAAa26x9OdwB7c+Qo1DvCV7TIs7rhnlhZ5ILLe1Wc+
oc4LZZ55UdPgG3rZLg3xTfysgweBH7X27ii61ubYBxg5ME0DfNe3zPDdNcbiPccL6KqAyTLrxItd
4+h+LxQg+5aA3YrjXO8POLibVVxEZjV3lK+5P/4Hv1R7qiSs/bHhWis1Th9wC4KuWmTkEiXRQnK3
2epzmikOEapx9oXRtIdPM55cm7FtKeQ6cohud+ZCNznAGPFEd63TACGhbATf7/S6nywj4tvaDTHX
V98aZchyblIQ/y4Y4ekY4XDp2aI3wmraduv3642hJzL8+SOSuZoICNhGIKyKnYBfsNXO7xoxMFJi
4wKe5/UHBBPou96CLSsbsG0OsRvmmGiBKMLmHi3CsoPtjyoNa/O2Ewk9Bkxzj7Ejy6jb7gjtjGAb
iFfu84iQBY1IcHifJSmsrutKFLccefhRaiO5xFOE8wMQMQWs13/ej5jtdQR/qdSJGZE6QoktYDGI
fDhcGNtjz1WtWPLvB9+toCuKg3hrdS7U4FtUWlWwMOaoKU9Hwx7y5wM0/E3svzKNKPwhmDwuIJPB
ayZFzbuG/o3vuRdFsTFS1idU3xLKRmD+riww0rzzLtCUYelI7DNS+0UCfKOSDF4T+Q6P5ENSfyBa
MqGkgTX9FckA9Umwle/hysQK5PwD0DNZEJ3njvk4hbyrqqNKWUHnddLISmdg3MN+iRe1KExj8Nf7
21Q4vpgUTxo4WDyBvj/kajpDeqeM+KoZxdmyv46JgmYDfnZkxXH7C5TX4Gdjax42V9AZfCWaWIYx
V0cCoMMg6RXxYLlFwLxGr6wIGawglzLdDVF236AwWkcFt/DfRHFK4hXl6PPAP5XCwShopFqBDntB
Myxta1dE10p+DOw0rEL6ttJRl19BNIY4+P46OhqF/2+iB7KnMr8tpmks2IlTUndLrnIhTgD/Brtp
NLoidxypNQ9W1fp1CmZ7I2pJbW7BnEJ3NDW1wYMOd5GW9dbMkucx/BtJpcoDbqmd9DYIgIGqXHcx
erA5+QHdu9UaDJYh4V+PHeHb24NH8EPV3Sr+HUmxTo8KNmF+ShS5NpNMDB78XccDLUap0mxadhLS
af1wM0RfQDJ3YSggncin12aPaWcH+lN8eg4O88cDoXF2mPsxLB8dV9rdFSZi09EzeMcnPdx0jz2P
lFspEAqq+hj0s6tXZ4I9lSzhrZnDLLuOk28nEoMo82C+uPvabNSptIKp0Bki06pyi2aTf9p24HVM
YhjUSJVKBTlXT7kVWMESz1tND3CdBroMCYuXTkcdRwVxiOMXefjUDFB9L+lG81EAdqTSiANPf7zT
vQfeBJuLY68ncgf2WAXe2TdzfbmUTlbzu6BuvEgGe0VH5j9UJb6pGxaDwJwf++JB/IkW2h5YmWeO
jOurPYqmHYN0KN54wsISQ1uGv7LH3LOOCKMv/A+SqDVZ2L6WoeCkBLmnRbJOvKgtWX33xQU3gSGJ
Uw7w8TQdp0CrDYNd5+KRDy25HwJVCsOTxistdGf+80w2txNlAXGBHHaiAyFrsJN8vKovzVB3N457
q6Oe46wPdVPQhDeJ6nD4Y5BX+VOiOMYvVa728BohlEK70nGH4sppRVk2fcnRYSbWHx3yBTmBxtKX
zVidFd7MsawQatigw/5U4dXOOzBGQ66VuTjHHbcm44eAWaNPFUUlQPgCh+cYxs1ShMHt/aUVjwL+
uPCQKssbuapOGgYfdQsSfdbpKmMLvvScWd5XSEAlaNUMYNW0low1FdrEicpi+fCsF9ciFbHVKpU8
3bHFKOmMoJGowBZB6iCgqy2KYM127oiDVtSJZ+nGx92v9G3b3IPfVUgg7tFmWLSlSfl6C2meFTKW
WeP8JNJ9aWWUhSTTWmMyOLVg3mfzXXBjotukOMHeIYtJu5sKI/2k/LM5fjDDUWQiA+QgcAZsffVL
TDW9zDtUEy8pYEJDzpDU0UwXTuXwXI5QxE0uJobeZlV8LSf5RHNMrq8kWC0QkQry/c5lLYSRtz59
K//SWSF68VmA34Wb79sL8DtBXlX7iJIGTpH3pO0NH44iDIm8WgqN/nPJGFiDdTCFUuS62Z8pinK0
5RjhwSV7d/cC9w+8acdobNXIECd+HMYT4VDQEmJ7Iqgxhskj5F4ZUIZFAvuCs0j0rhNw5awxIniH
60HaNTKMThgJDCAMkoAX9COrptmZUqI8WwCz9QSt3Hx2cI52ciftPqfp8zuZ9OCt2Bs2X0QS+rPZ
TBR6rh10GCwwS1E7UD/M20Pw1WnXA1gWpwtn2YeaIGsQBsKkiIYt73/9gd0/HBhv0XBtm2VIDXUJ
SlVg/DDTdNOUF7ZMAfQTwaTT9VsaapRBepo6Dd3lc8p2idDhOpjq2AGgZ7TCVj6hzdgi+5B57PT3
I2U9LtRXRR5KwBvZISm0C8hyUW0yXryIHNE7ozQ2bQ+6/CHqoAC2OgtUYjtmKR3eM4PYTregvGIJ
lnwjOSE7vvreQYmd1TxZCdHA1sBsW9hXpy/T1JJ+qq5yPLUshdxhzNLlqKi88Bkpa9FVA0k0IDFw
+056dzDOu9G+Rg83KekYrN1KqWeMCyGo74JfCmCIJXDOaUg8ipDL5wzMfz7AZhJ9CGqIYqfU9hTz
qJcKsf6XKQcPYCOf0ufxBt9I98n5L2gYMd0pc3bjex7o1EccUL2YbFeqf2VrGEc2ZogNIB9PVIvu
5gE1aY3aovrWFwGBL87sU2MiT4nRdP9cTobsQ6bar7KLUuc6wpeb1976aBP0rv4sVwJux2oyaMMt
QVh6qb072z0KwxY8dzF4dGFza5fNiJS5saXdaNJyxT9gaELvNrSXLI3NVWUbXJMmzCs5YYS5bMaf
wA9vr68BuHInZ2qxajDjYCU5eqQ0+lYCXqw4opBYTT1RuLsSa25Qm11o0d44TggzcyONItAU+CQj
1IVapcm+DW5HcvjBKNX5+rwTQ6v00oKNevgQ2p4XcLWECLoK8ExDfVnq6g3isnrKEsxXSBdmQyZE
mjFPvtig+BgMckGnSa9alKUGJa1dmKKgbgHpmc+7TMLWS7A/sjlwEr1O1k44Ns5V54291AGFzK7N
hNxkJwJHEpymHBQBKjKmswNplkdWnFOcETtffj/3m6ID8Dvflc3ztu1DcvTJ2YF58QMBUzH2jsDu
O/vx2kHd6Ryod45mG+1nh44yCTg2iJOgHCa4z2ICBHodkLRinuAwhcg6JlAksrTXpC8X8el+5gZv
Hxes0crfcdfiMoyUeAUgAjISZA+smyF2Ix0nH8uHts2PvCLjTwUF35WX+DQNw72KPXi6atpRVVFk
1MiQksZfwrloY6pitg1kBdDd2UURvbzTeQJPpharkcgTHE2g6D8Lsb3vxRBZduEXKyXBkS2vtxMC
/5C5Ka+s3hlbOF6e+38JVCq4ZteA2WYqEZ5902zfKkClETyQzMvalMUPXxzfFCppGQGG/VXbAppG
ScTAzbahkZOjp4/aYrFnAtT81v+L/mKopEJy9jILFuy3Wngp2lYi3uL4xiU+mcfOU9HSxCAetFQE
4Rc2c/7FA1y7OJkyYwV7esX+8f9EVdv46BWEJm24ZnkXPcYlnScnghvOnywcjE8vuVIJGDHHo/Fd
cAfbI/E9NsvXwrFoloDt4xLGsqkYNvZ4q/Tp4yTgjBdcR0v6SurXlT/0JxBaKbqNrOZjuvLmw2zv
2pKDDtKyMh87rni77lF35W3SE4Sh+9iu5vCZuTrIiGbwTeXT8im/lpbEdXFxOR0J5ShMexVo9qtP
rsqcnbinrm4H/eRofmyZs2VU6drbP52CFOp8HgJHQ02K5sjIkKvfaioqU5p01wIqvA2K4v4+/mah
baORDTHcs/vvW/jnxUMxLc+HD/ix9T86bp/clCRYs46IJY1YtvUGE/NJgtx08UnpoV1bOD+IKhfK
BmcUUexYnvPcNZR5GFjws23w2J4k8jBW2mcejx1rw5e7cvWCuInJKDwUFhUSwmavhImQqQo26N7C
E+Xlg7lXAQzqr9NVAfLCZGzRl8paD38IPlQSVc0T7l+a3lfhnG4eeEUnaRR6VXxvW9E/B7N19Plr
tRJhvZ1zAewf897MilETmNZeJ4kK5mYoPPQ4eHI8RVoJUgtDUfXscsUxgsDjUgDfEcCXi0fhTMRa
3B5F0YSedcdVZCXMFhc5u4PmgIu1DFv4dDbD8yWR4QOJxwCeVwtENlrAirQGE6faPgVt34udqFSo
0vxuqNuzWkz4Kgx4LHjYd2Fgc+gTWC745M24LnG34JNdXCFQZXoUpQeJonKQ9Rt41BGUyHuLD+Bx
qTPb8PtXFKNbM1ey5kLZyHr2R4lwR3IeA3AhIZrbkZNbyMAhrZ3qAV8z0z5sFSm5MwgXabPf+zPu
UT1Fsyg+0gwNIFSlF4AQi+b9lvzl+KxhtHY/tSKUOWqaYQ5ZiiF5nVJuIFuR0Uj9xEilr2KtGBR7
kCOKUwwENHmQ3IAX4pqvWqDgnFbLEMF77MDSMGfAFOWsGtgAMwb7vOj/1qxRBGVhG4lNjsxBdwpG
u72eJqJVZ5zi2VYpcChkiPt28NSfmYUuqNyEoZZABavIBry6ZAQqePAc2Tb3p9whQRjANX9apcOe
oipgPnW8BU3DjS0P9Rv4hVVBekm07iBpjZtotIex92VKAAoCjnspKBDFJzGiCiY0WKsf8z+9ejfQ
77sagKN6bJIx+wpm2sB1LiG5cNfLZbnIoa/EKLsII2/4kMpxzP7/FTP0uHE9u6oO2a9tOtlZ/hCG
M0rQlWLq3d3DLVpDUN6Kkr8zrpWoAuNJXr20KTDeB6aS7JLIeDDZ49CcG+diGTWCs2bpD2Dxio4l
IEJTWKX3iox2WOPJVs3U6xikIKFlpvCDpkAdjHTWZ//suKn+cZp3U0mCe9jna3V17AEUkQUVqnfi
70vqSHbMY2fKjjPpQjH10hu2oQL/xUh8XET27eKSk4THyiGqNMbtGGYQUQw2xDDID2mzQJLuLhAo
ZWrMAhm0nLuHUlp3TmFrzAi+F0IMNxQRBvlKoPydu/m2HNAgXkbtWUepWO7OqFimPGFsdzojVJ3Z
omoK8nibGZKajpe0X+MOlYbRkoHUywa/HiWkyJImHEMFLRrB5akEIN3AiQh6u/mOwtU0p4B4ry3W
mhiU8L8g3L8DXkrlS/ecG4wI7Ez3d9lLzfHQXcUGxMVl4KPCnuDImX9KB39LTXioOizorOgR6W+l
+a4s2gaweSbSy+N9dPnXZlvZ3wCIbRsXwyJnYgDl7TeP5Onc3T4vOq498avFDSy6g06w4UQHAMob
xhkNNTRxof+cKWOrUw6091kXrIJdz2h7jMiQCh1Etb8VahTf85EHoPz3PBcf9nZ2NWiwuhjlkSIg
XIaBT5/Epv1stf/b7h2otup+neGpGfh/y8n2/XmecnbzrMT//ZOsPXpHuNWQLGsK/JdYRYBUokcg
tOD/bFIXm6NHNzdd0l7sQxjvz2VcJBty7G5od+899HY/3qIaFsJulSTCaufOMdb5wXTB4QBdk08m
H9TJiNS0pzeIkRoOicdYeSQGzwOrbk8mmeOCv5m+XYGTpmM2a14YLzy/xl3/DGMwWOWubKNRtQWS
o+CwiQovc1MCd1uF2zo4q0VhOyHGSlGBdWuPCXH30lJxs6YjXY5FL5Y3Us+0P6SOnZ+SeiaVNLPG
RgFqGAoZYYfkWSEXEjNkTI4LEbkVsoqHQ2SAeBLedznh4iPRRXWeF/G8hFKZvBBjeR2sljLQmV1I
Zp/oxGdYCDpnMRb1U2CnmnEVAYCCvhlCBce+9wfYJDotIGuRs0hroWYD5E0dFrJgizdXp3TVeJTi
xH2MiPXPgCI1MM2h9RX5fldYggKmJStlS/GczT1JJVlZUUk4xXseRKWT5mbgRoYQOW1opWUjaLoT
P0o25JVVlJaLr3WbGdmeIQJSy94drI0VoBoeicIBgYNRu3G3gDuRo/4SLY8rmUBHSgMXvG4ly7Xe
2mmJk3P6KG2Eg7ABcbt00wfZfhd79ujFelPvSRI1QNrqf0Y+21I5FeWiYSqfmia7cfRNJaKGWE8d
nxsOELv//eSUi9/oXHaMnpy8trMq/uQkaIZkYOFl33PwpIZyamOgIY/YFj6GVJriT+EzCyPUsAHE
uGkdann5thekKxHLwHpqFYzpOoU+FUjb6i6dCzS2Uhi2NWksWHvQSTCw5dVBjAeHESuKyn5Bfnct
W3U5fu2usHA39UVQtqzhMzMlXl61+m0+lkb2UpyuhRhNhngnXuKEbpHKcfkbaiI7yaLMMXrLPZ3D
GUK6bnrKFLcJp/SXLcBZFqDdmR43TynFSdGBxVqtXEPCkHjxD4wpIruDlmSN6Mno9vPxVM0+iuYl
ydRq7NY/uAz2jYW4VsdwbeykxaYvVDqWUxdyGFNPh6VSp5OIewc+9CFK/E/uiUZZD6CvfNq5NhTP
MtqThM5CeXu3udiS5GSQKVErm8V54Dz3ZtMHLkDcLkAAhGDvo5KPEZ5/k8fP9VLUbgRAj3vwkLAk
zxBuHF43JdNx5zH9HzSNOQu/4SXymBJc5evqRT/5hXnKv0McKRM4PRA9Tf4W26f1P8PBToxrfB4x
n4iNN3BSQi7n7xH2V1gorVOYnWI2Xdz1Jek8RaDPm+b6miYUq8eSG/qsQwZg2ymnvyRDdH7r4Puo
aS8TtrrFLlYATZqYFmOsQgSYWu5FDMJn+Qc8wJyGuAbPac+vUtVzZfSVXWJGH6IrcyGIiy5SzpBe
Fr+qTUlA+6tWops+CDzLEeyqGhoYlAzVtHneTjkZU0BkQIUoKGDj43S+A6bf5Ox6lJmGUWzexQVr
k81vL3+qXJhp0vdnM5tx4rMM3HywZ9nD+VuXx/MA/yg+6EwheqPMuvq12Yj2moKXImxnkRAuTAU/
p0Q85FUd89uLg5NgGvyEem6XpQ485pHrKpTzTWHCywvI8CCFbqo7JroFJN4IAB7xXFgjRw41atN1
Ggg06k7dEBGeBvsYZX/QhmbRcl57MsEjbc3XRzezz8pbxZbtjrWpd+6wg6uv/lTbS3CJF9H/Ww8M
GBmBXpkKb3I25o3nVZMDoTY8PT9PKD3jD6gF4St0dGQJTLZYNyUa6TWAPopXUP5P8TPzV73KqPkL
qd5McFCxM9vyZWzUD1S39GHuIoij8eJcXbaqdGiPI+016AoClZTdv/t++zwrgvQeOFzMSefjJSS0
L59LiB4LCuPkqaG4subxQ0QnJTnTIglOnrQ2vaCaZY0LgJjROYJUNFeZUWxB68ewqdBJHZZGUdZL
Zt23Zkz9RSxs9lyka6l4Dn+PRZrdcSISzU2sra27Eh3y1sJHgkLJCZ18iVvneWmnQ5gQ4LsiEqW2
2C2Lrb6TWSaeQ5bYEWnl2gJ/dVil7n++WU8KTUtf2D2zgFbw5LYJPKBsC5dOjGuRlGG6Q27crhLI
0OoooIIaoae/OGelxW20k1uIHZn6bqavrw9nMwysrLQn2RTv/JbAGSBWL2XpMY0fQV/sFl2ke5s7
VEcWpCoFSPge2Qq9FlJZF4ZIBOjHpUhU5P9z+Rgr4Z8kt2SI3vKJ87+1HoaB/hnGYe2z+mb3+cc0
xG8rE9diZ7qltgCXWLYxAeEbV7/dfjAMhgbH0Lz4UP1InimftTqRRvMBJ469GeMiuBmLvs3WzOHw
BJF+gZgtG8kgi9m00C7dbvokd8QN+23j5Km5hXWjakPGGjlV7bQLmWZN3JnmbhPJz3ghsPNoheRE
yxykvb8KFn6VnYnpCOVyc1Yim0UNaVOj04qDdry8o7ejAIpN/ZHE2mqIB6qkYQP18S83Uhg++ubo
hKKcsfUUjl12l8Fpfu4V2e5U3XcNnLLhnyVwG2iWwPjEZXgcfMcj6eV3Wj3UkPlc2ZhN40BstyAN
6Uv223fdXbgOYvKx8cs2msyRHTPRnIA/Al53Vc7rv/nmkkynlbIZar1P7J13OfAgvkllC6Dd0Pjx
nSg2KB9sfQ6G7ID7qloHuLvO7bdGb/DeNfYcndSFr1cOeiMThyXN2eGwT9/j5r6gm/FJIT3uoJmw
4GR1YXuiMZ29I1ZQmGGKUJJKxmJ9b8VhJxiNfmXEeIP5WePEWqTeUljSg/o+63bz9wxvu98y5td6
PBPjjY/gi1HK0wde/3+6jyyXhDZmNq66fY1YZi/nRsUoridsuTg3GAUFjO2ODzkEFI2/IVzo9UFA
lGhbE93yaOuKEGeNAVKUG/mLqkK5+K+G5X7Fnd6F+YsJIDZOU9exLPb12Br+ZYT5opPMYFyjTcE/
C3/XkULsHzVTK+QnnYA+NcKd33i8ElWZORhCeAtno6keY0pSOs0wxKqFbDtAEVX9HJd2irVb0Ap9
BcTym8tA2BhiE0S1cddNh2/FsMSsUyaW9I41qKFRNfk5HQ0mlTCvMoLFhUBFahriV61h2POat2Ai
LcEq2fNgBPieuR0ax255eiJ4xH6bRBqvQrfykkzANQOBR2zHIHayI9fWQ57JVLYYQheZmJJT1upc
tkjAnBQTXYivwrJj9D4RwkhpkzMH97auGbczh/Suygg9YbEZTMZjKvo85GNHUo9vLdYAisJzbtgR
rnMnyRwER2oEQiASkFGZS4QyEotGpwXc+gi/xOIjwn5BNdn7vtBRbcbVgaVzJvDOxOn62pnfSR9H
HKpFeYixBU0THx5+XV80fbrkxX86zFdhhhpK04xRXK6AU69h+k0ta4LhQ0P1L9xHGdA/6jbcCPwj
vHZy+ci2HxMXcqB9DSNc0eQrVpBh6H10xNUq9WPgR/maFpuMwmpPfwADOO4VWTmGYMXJ82RI59yc
YKqaCcqsRMCXBV5qTA8btB5iA50EHT5lapEMZwxz7ZwPmuqgc26FCgYg2z0hM39l02dY6SG7vVxM
P1KAVDFCjcDWhuebGQq0yb529BSEVg0dv+vTWG7HCkLPVaVP3Uv5EAjwUcU8AAAnYhsafNZPy47s
JZlHM/j4+RWrgx+JKijq5JZIE5cMEzur6tiyDNDoQkEhIiewzJ4aRsCh1B5E4uduFI52QfCnMY0u
321z2qbzkeEBVSlSSum92Wfllt9JXdw2dqnvVF8pxFpM5rGoLRTFqUrQ6dogDNhrMUB2MFRS4ndY
vUXc55GIhQd0DF8D5FvSSCVBCdGfQaG2H7S6f5soOY+mvd4Ziaj13heVhV1HtZJBVm6ZoqaQMiO1
9znTpBzP8n0sCeRmt2dubKxdI/4NrAnndiMrIyYc0qkuIBLR8/HJh12YiGKa8vb7OL85HafABTVA
tKaZ47eSGvD07Mp8D5/47XiHG+kSQX0/13xHgTgiKs/uXAaukEDM1WHeus7mPCEc58JeCsMEuHlV
lEdB1AQPjkk/MxazwMkXnS6fFNoBPUBnKPjBeQq4PmQeinYe6AP7eDKifXaZwjUW4IuwzbvTWOII
lnf6MBGwifV1ehqOAbNW+KpD2+qgXPSAKkKe7GLwAkYnoF+pH4dRAr0+V7JAVfDVl2pvrv52lX4F
bMxC20CfJeLHJKLKS4Dky03OVkqL11/bATmPS2oBQmc4DOJErUJ5LJhpDNF8YKx7VMG513dOXO/N
Uhm1uCaXU6Njmr5719XadDxhj8gZUVH9naP/IlNvpIvLOBVCSRY1lQi//ZZRinSxwl7Ils86N1/f
Xawr3q5hAMQrLQ7wrg/K4PocZTriJzBn+wc8taZX0GSygZLb41i9octpId6CDSkGTRLjepR3aaCp
M6cUJyX1oTqIzfSgGubmGzp9MK9dw3GuH4CyJr7sYefIcZ0hqQoB5a3oqIDROcAHuALd7uVhp0XE
d3Q0JfTs4i5Y6PePU/OF/mnoAadz0rgTiDJw3lDOwIORik0JF1U+Glzr+u7gP6oChMh+p8RYXR3d
TXNIEnUGYww5aiNEYhM5Rvu76CNG9rRmSRCaM+49pXMvQJh7q1H2rAGtppI9H/hP7rlx9s1UoWIU
umYaopwYMmzD1cnIv88MJAGvk4ZG6xgmky/RZ6/nu7BCohPhd6RZKkAKGN+1w34m4g0MLKQVGVet
rnvnyt+iU4Ch0Cy1EYEVWbH7j1IaSG1zu1lIzo5SG8NFzgkMEZabV0F6pgXXowMdqnrl6lo4HTCq
Wf/wG/VrMgF1jN/65N1ykGRPi04ed/bIp5r8X9PNbJndVrJWGNOsvO5dzD27QHtzX2lhUJrglzFs
kKs+lBHr1aX9Vm7fE6Fme0VYHeKF3XiQ7+K/cUKcV1CvyWvHmeLSs4vGX35CaqTMy7hBAcIK2pd1
jK9b5HGlZDhneXwwsvg8ZfCt4loYQwTa7DDchakH2PeTN56hHibltFL3K4SMd6Nmr30jUVUmAtAd
GigS7y+XmlQAuWyuWma/3+3ezrGgDBunp/8OOk2QsKRwqhZFAQMsOPEsjcdbqeT04HjI570JJkr0
qbVoLeIdD3eZsFyDD0v38i0K8wpZb5Hv3Nv0jeDE2ZFJ2rT/ChYc2AtBlMcV6c9yC91Ekg82unzJ
gmobg8D2Ngv1fWppjK+/Uj7qFEXzYSMGep4nh+O3xHMISGAX4NUHz/YfRG3HChIsoCui+xJZbeI6
r3aW6aEdBAAjOmN1hRDBDTBl6+/RCz+qCZSE9Wsg9dGSemvklPxB94MzpaHT6v08q4D/11SMjdiZ
eC+3UhLLDfMeujuwq1NYoKUF5DHzcPeS2iJjUR+KUcu8Nb+LGG3qeAPvzRUNrOwVb1Q3bChK470c
is2Cxpx7wfYdHlLGWZQf50qELCjRKTqXMnfr+NbIPw0DfLIL//RsOjB2S7iH9P+LSzJDbnw2u3r+
4dDH02iKjszaX5URmGW9WkrPYvwLu0wyDm0lRVXid2AMcrUrqUqbEI27RoYBb7o06uet1gPFL8/A
SvSZ1kaxIsbgZZ8afKkyvYO3SfTokmZ3gLrWaWBCcL0AZjgW96MYMeW1zgeuY+Ex9VV6EauMOlxB
RtMmIn3n9a6bRyR7OtuTX94t5EnxOigwhyr7cnmBVNw9ra9JP/9Ytc6fI4IVbItLUgk+2Bh1ACxI
5YDGcdFzo/dWuaBFUhMzN9kuc5eYR6fRVJcGNAA3WY7QLVzsq+3UOuRyLzN8ybL2o7kWtcGcl5uU
8TkZAvqTS3lzjCeGgGHJpf9Z69f34/KtbLhGLhe+I2aj6k51FK/OpThkulue9CHsuFm9bduBg7yz
OHCd5xSL7okCRYtMvdbcuQIqwfzyLR/tEKP0qOhLL32uW+sbF4YtiTq5RVo5vAufh/7bLN+6dtjl
3syIUnDQlgcgUrRDoYJFomRPlrWbpyi5IOJrrV0aaJ52qnqPI1GcFYYNylTFDgfXBopafda1gPjy
G6W8Hmmzr4JoIH6PvJfR/T3Tj4GM8BKwx3lw9EBJ9ZC3GhawjuQib7MIaekMOBDQhdWBNmxCErZL
MFhLgk3fjcDSzTG5pX1HGga+e1CxU/S67BCDuF9nv5FAELrLgSN7KKQdXWFBKHaMTTsMgs7G9LV2
noZ4GuZRIUo6QNAc0lUO0vd0jXZI5UrAEvU7B0wXx5XhwOZkwI1ZnKQTcJjjRxrkInPB4Ar97CRw
f74NQ4LE7N9DxR60SPE9897QQdc6K471+V7q08HahjecFybnbDxmVoOokh6K3wVUr7blEXqBA+iZ
+I8DUDZnQ7I5ILtK3FDaPjV0o+v4uPwbUh+3jLC6TnGcGwxJ4A9l5CqY0NA7rb0ndzpZW0ZPtrtt
bs9cznCSTVPZSDX8cWX6TvntDMf8oA8dpjuiwQ6SzC48uNVSvY8SuPVuSqzKbC3WE8k96CdWdxWd
hUN8IGndD2G/zvTzWvlAliowrn7Zl3qifbuQ/LiQ/dd1h11zG33AQIObr2ZBYQzEmLlgebZ60djU
WiCLPFar8mjp8kdMHLE+6Rp6YuSzAIfm7JQ+LAO+ZkxQfCDfG6ZlhzqWqoRWO/elBdGAko3SJQYk
oyWFKk44VoA2Z1UnaMTvNmVJJYDv9OT9FrHvALqdq44U2brnvS1S0jfj7wCovU8iSCcYSFGiyFqn
IfZCV6iyseo6enoC4Evrj4krNx1Y7lYO1jLkOO19nHeLmaIDdwyk5uQkron/0F6+/mHEztcgI5HV
1scqrDjELnYaNNucSBR4pgVWncCEc6J9aTMTHd9sdkXo0Rin+f+Z8OwOjpjswRglljhYwe2/3zWa
2//rBFrS8RE1zYtEKBFcgd0pMiPZ4V4E7lWbGWHrc+RwtA5FrlPtc3+KF6Z+mUwfnvVEzFA6CN+V
cLtbpDlfawcYJs3vc8zKjegMmOHmm1M/P3nzvqy2Ra5jXH/QHFe/AQHfAnytOkxPvZ4X/CGwszr6
E6bTVCvmxKRquK0zMAlVJq2jTWZQGuCkoVfpMK1l52NRJjpAk1VXSM8IcatSUifvjn5xjb9XWTB5
iZAg4I+YT8sEIO0IY+hA7Bq+R99+tKzf9XRtzJno4prAqX+28jlcXgg5sim9fd5cRQwfFhRP8V3Z
itWix1TzLmX/f2ZmxyrBm3zkdoDh5FWuNyzsWyZiqhR2te6IPGtczRIXgzz6pLHIKef+BbuezWsO
e9aKI4Aa0/aljVoWfeJK11WNIa98Z4f6jtWsv25e2chW30uwu3YY27ge3PXvu71+vEw0A8Wqus50
/qLL7LAT1eKxuqQ1143eIIEvXoIZgpKPVyboXEI6J5nedVS73As+vCSCUqd5/bGBRIydwdKn/FNJ
vfF9vA/g+yC0ORlWC8kKQ2nv9rnMVsYlsGPjiVOTVQNfL/S6uDTYnFmRB89OsIGudvyMF4Xm98fL
yC9QG9sNL3mV0NeAgbphCK82F9VRe56H3e1V//Vh5Lyu4NLBTJdlJLAidRqI29os1jRY2AO4opAl
xlGzoFYRbRWUQkp03FyBLKOe2f7O0nSKcdOCNpO3L3ELkKIZeuwRZ750iIVtoCoc0/sX2f2iMwD+
iAjMvwK/YOjlmDxl+jOYGBojOqYfUW9NMiyZi+2N6zdI6T8tWsZVOkl3lf2cothzY2hQVIm6QVTF
DeMO8YdLEfa2eZ4XRh8w31e+IgSQIWs4Tiy/FwgbufZJi1bc66I0DJvk0xDL68KDMYhMCCIMuBVt
82QJLX0pXYu/mWULZoOQRCMx8OA4Y8+k9ILIInzSXwBcXCOt8BNrGE/egvr/VLqT5SsxauOuGBC3
0E4kCiBLfIGUNMNX/K4Wq3mbnZ5OdDH1N8gIDxGv2oDIBdrb9n8ySe7BjeHMS7OqyVd4jX1EzNCL
niCEsQs+oPFPfDXsQAhqsCcnU3H0LWSoNWni78QzTIwqBbRN97tPmitAsAwUTTgmaOQfRYwJa+IG
TXj9ZOMK3UFc/ETiOotcPzkQdcfzQJIGuCwGeDNVxNZcch9g9/UujbxPzW9vnPNWcp4vK9iHo/Ab
mgAMbtwyLQxKj5tbtoMX8lDdvx+yhI/QilMGbNE9XIVfUsmtoJ7Zl2WvugYDpd2ZmrrAtUFxCaeL
LFAdtlUIh4iTdc3jcXM4AXT3s+ATD9Zr14wzhg7ZL5ZNm+OrOkGAliU/Nq5z0xpxRHQQs2+uddCn
6DOC1q3ETmQtfO6TneXbCYDEtFGK+nnenHaSZ9y+eXMpa84VGblYobg/ujjBhaGcQ1CuKQ3k0hPa
HEJOjyT0N+GlTE48RlHuHht7241meyEm0wUfEwX2sgwE0ZenT6drmBg/X7Nuf3S26IUBlXgGDJME
Zp7qO8DVkGmJLk1QaNndgPk73yYF8s7usZ6udy1FAj14zMjWeNKAZ1ojJqr+6b6w1LvbciTe2yUg
uAlS5G1pN9g6dAUDzTnxj5ZFFhQsUjJ1JwAHuUuFXD7TBqqDDoe7ZeyEhD3fCH8+wlLCCxiMQluw
rSTmSD5dFPuAFmE+mG00Q3R2Rm3EyyYyHONErCoLWAdn/PW5wnFEliAUrHDa1+5/kO1L+2ZrMQg3
0egEEuzlOkcN6JemUohWCqxzyf9OwVSXR5SJ9Psh2LTur6uZSjroLYJWwvsfuuHdg8fmslsa6Del
xGscoYkZ/rp0pZaPZKNbVGZTdHAxpYebD25rWJ4b0+rmLwZDrosR1aI/5RaH6/6GH0uHuPl618pF
0j56sfw9pvYv5E5pj/FYdZO3o68iyx9Jz891PylMQDkg5VhjxOzQ7XkrU/qK5FQiueWPgQr6zZgl
cqLIFT5KBzzHf7ATBnf7COtud40SsoOg92foqT3BZkZgugFUDgdLU9y7CmlG7Jb9E+IYZf8Ipt1g
G0ZTCUpd4ds0xm2WNQZWXeOVfEbIZ02eGvdOmY+/GjLTDISc8ZKjQzKjZbrCcIToO25HuKIQfwGH
j83nRM06XuyrxnPRcWopHwr/OtFtmCgyxLawaqp1KUc0Qh1XMbJtrlIRMCMUyT3yJurd4qlmL6wP
GTtm7yJFTvRKUC777pzQ6TX/Xs+yNVLW8zBjUuKMONSBKpYMaB7eZ0Ecow6T/zqqbusiSdAXgAiI
Vy+YKqxafGNXd9mIkcCVx7HPGG9N/gnakRJ5pOTHxMce1oaet3rVjteUDbAzdGQRqMiO9JCDMRwN
mcXp5mb4KQQI2VkDa51laSE2wSjb23jG/O0DS58xFI2TJHvA8bvRJII1KS252Fx82C+Lnotqostb
520wB4A27mUISkPnJEx7/ofXkhoiB61tsBIQS5tiZY5s/ikY+d6THNuhdZuTMXBr6DVjx4oDdSf3
GD1ISZ/iBjm05fsxabWlFfv8CH+9FPcE43P1m8Q9XVjbm7RNnqPv7lzAaFYX41WAh/RzyY7UpWUa
iglZrBKjLNpsIMI3IwlEsNpicUh6pX3KivjGE4P10b9rQTGcBEnAQqOmvuYwPMC5tbV3IJm9TzUb
ezVPGsUwYLbEIAdG5bAisaYYpYb9ZEMcH0Tc+PgeFePlI3cLqLbRswPTICzxBkpWWr8i13hHuErP
KIIqiXp0iUcWltStOOLLSbLW1tge/zqBFVwQmbss3Qofi45MP6S/yqkwZ7347EEAj3tHHNLa7pcw
JO6R3CG7ocH9JzSVfKkZMCDoiKsLkdXzfT0PKpn4VvyU8RU6N7G4YMKa3EQ837Bc1jTouQUp8U55
Mw08+KLWfXzuYmLexhVOpz/1ckkqO/ZjGhbmr+FdIBOVuf1QW9oHdc0VvgfG95WTnnsTzKWDjqym
ojMe6rOjiky2IM2z7GMc1IuLdigq0B64ySgjAEr8SnFCnUjrEw9PY37TQIRdTNh0zyn5FXHOeNqD
eOp/AN4AExJMxggX9Gv/mFYyptqqTnLyeEWoTSYRsvIOvz3tiyEzDVerHtTVDPaCnZqZ6ZGHaomh
D+1oL8bLXWsXPV5EmvxFlJZY+a8X+JIdxMprTk7I/R+ZimYEALlqEPjRIE2e73Ma5SIyGPAQjoEf
HxCtryoiU9bTylf3gTT5uzrBYPmqTcN+RXCDUAGd7vIv79JRd1lKHMMNY6uUbPr+3fOrDWNyV0m3
KcFk/yTYii3o8F/Xdex15mD4GluibKks8B2R3LHEWgq47nplqBYgTi0SfG0tq5rn2tP4GubXcRfz
jxXx1v2+OFeBReG6D2BbaAnXDGd6igTEIRojV0sz9VUKTtqf3nrZtYbwusDQvAVgpKoxUMWQ08hd
icIzHbP2SghUPsNUuSpUv7KGSXNG+0bEKGm9WQTTTQ71ZIz50Fbc7WZVV5F4dxUQBtzNJn2V4wsP
oxuz0YAzs+hjlBnV5OaLzmbBEFp+/sDWAxnbfVKPyS/71a3Fnd5H8TSqNZy67hcJ48zkxeZhIFIL
PW9NBEjzsG8OZEpKmH8wOJlohoyB1Z9SmV2g1287TTqKPXkjIxIOMw9EgGr5mdPsYRRwcDRfdsFS
1syr3gprjyfsXw62X2muzVdmuSjKMeePUWXy/VUQavG/5WYRaWFDssWCsdsdGKaP9FncNlpk/qqP
WdyfNjek7PVNNmKVH+DJ2AwWSTrlKgkh6OHnZY8MUj5evZDAdhTsOvVHroV8Hu/hhcWndfynzvWZ
5l1/o0goZWxernR3bw4ru58G01AMPGdxXCE4n4601A1dM5OBoVc70xox6BC/0dzCPz7L1cX4DbCX
h5fd3oUyqIU/phG9pg8GzWDyH/RkYhTQwV2kXKcf52RqFNnJ7jDwys9vhR0f3W9gfNAYsYdnLd6a
bY6Gg4OdTJMOP/8EUQXWT2m9MC/FPOYwMhzD59M7YwXxQN8S+EdHJHBhr0KikwJLCVrsESih/Teo
mzSS2qjH9CnoeysSTxedPqS3CVDrZuS4q+Oj+nbpJQm+jjSCqOT9VgW9agioO0rotPmTiHkgSIw5
3C5hBTo940aZxHvPlBy8PSYQPb7Rnvko4Tw3GzxOCDVo2VN+cA7EeXFtrPF+ZQGFxuLMsAxaxFq3
Yosf0Ac/wcoelQkDsT/y82NBONJpdKFpwDj64UPty6pTBLSGAfPQKeUhhzc6yo2MTCPEYPDIKl6Q
qAXppZikwItqnWmI1GfKX4pASQU1HncDf6usvv95OShmz4EPTxXkb9+ua1vqcWl8jddtX32baMXn
UVI6OzLwrY2wRnR9105e2p2KLskrV2kT6l6ugqpysgyZeG6o3lP0Vvsl3oMTS9pWIzlwRKUZYTxu
iPNWKFmvIv7gylcnSgqMgGUBsGnr7/UF3FByoXNrx5lLxBtMlB/d+VTuPZr9Ul/bwMjus4yKPCg8
W0tgVbz9AFlZEGRCvMZQjbfE782ZJQ0mTgdJ5NlqVK7aWexOtS8chqiYtK974ABBSGyoxmikClzk
x6emkhb3Mai5Ot2dKMA8IQ7BG3lg3HOX0t+tgkAV+skgt811pMZ6zKc+FSDQlUL6IG21/0jDj1Ks
MvNYZEeQ0sixu2QgmOdJyiiwzmaROEtTxFxQ4k1Y7avK6RkS/r8wfd+rbAkP3v3CGtpwJTAkZZJg
mndjulS4Rf6kDMaCxjSc/sSjAoq5zUtkPnEYqtH99OmLUqnhokS+iBxtUBx/9H5DZ+VMybJfL3w+
J5CJun9ww+TYwhdYSPKDLiz5m+iKb5wdkbuXXi3tFbBKtSCCIWSVrqvh2HhyhwaqDvVV/vfEtRhN
W8O+nH7Z2qcK+qXXWtpfi+qkuFC90njYuIci0DC4MyMnib6neRHskpmFaRslmau+1vb3v10pVNQo
pkDOmevxaDoga7d6BZRTnNct9pLfgk0LbOU9nfebGTT45mOWhY+gwqeY7xX94ld/Rczm2dNyJBuU
h5+ioI4zmvuSWAzRHntSMn9Io1JnpUwHQnQtRyNiSLL7SWDOBTikS6C5xOxFKufy18GyJ2TwdjR+
tc+IuM1oyOXnlc+EfufFt9eeA7+jvrOgHfW2rjbrNPBcwb49zaRHVanbE/MwV2r3/XaN9vkpNk9s
SK8xmhBipsCn7ItFj77PCTjZhKFnB8noo1TP7tL5edwdmq3Ta0t/hBBL0ABQcBZBLpkISurC6yjA
Yfo0+UQMVDgyTsUWm8Gefmw6HuNYgBDw8YZhHzwfF/ce1D6kKTFH2+HwSgDt6RLmC7sC0F0Jj7EF
CTKg2YrCDu1fw7a4CjprPCY/hhgl3HITRWNsORDVqxlXZirju91xl8jozlUJ2EztAfQUAWR3A2rK
QlT82gKivWXj/DpkAje40J/9ve1AGdr1NCv1WHfGuSEuoIFNWkzHMUpdNKXAAKREbszNI3MyyAeG
sreSFkOgEGds6vOnnw5h6loATp/DYASecO4y3FbbFd+7aFJkSuw9vzjOJ1da59co+E72TPiWIzVQ
nJo1sUOeOF/RIN2rK7RSHnwBvBnhse9zb3C9M//pFcYASrjetFdEbJI4PpNRSEDuXnO5Hbir8FAd
GjhYSp7g070Da5jSTvQl6PVmm9JJX3b1+l+GNq9Quia6qEGgWONctWflXIi6/Kef5H9BdMfdFysW
5ttILUS2YUNXB/aDuoiaXmlVxddSQ1ZsRxZhdsC863cSn3AkKFrmaFgrtjAU7T1cQ+9Luv6+P8VD
Z270co6jzBxtmvOgofF9yhpTRlE5tZ4gaOEkXISURvFDpIOV0NI+ojfHaFpYKJjAAMIq6smYupua
e9GOtIfpenOudR9WEj3H3OFiv4L4c/bE+7/o+JUxf5af2GZ+z2k61/u1vl9l8OExo7lLts/6bYG6
V4mu/OGMKQdZo/K/0LjdYesBCAcZRL3CBNObfPxl7nYVUACi7qZpAl5L/l0s8h+e+wfCSe44cOqD
HX6ia4qsV1w/RQaDk25oxMfqal2mf1+aFSIFP3FtDT2EXCNj0ZNyHvz871ug4HWQ3NhefGAG8fNm
C8W+S5gDEsTz6x+oJauacyFu2a8WC3Crmi7tSGUMsc+fqW2bW7/NgkDDU2k1VKnhtMeXCr4DF95a
Wk86TEq6F9Xo8ucOSabLsGlpMFqBnQoeoftMnpsjZa1TzYIxqmlNqytW2IctafqxJBK177jwzdGP
m2VolMQv5QckjH0pho07sykdk6Iu1+7uyn9zMM8oJ3XPtAuTgXFUQ9Q41CYz1I3b3/6Uruae2jRW
uwWla6/EZcgMHAbKWVc7CggvsLTQIpiJUhLNARUG1j0ehfFSzkYrBGukvfK8e7c+tp33uWvjXLei
FlIFiFAoDG87OLFA/3/M5wNfWbUNRKTOHXB8t7kHt27T69ejEWb6agcOz+1SGr00X0ryR7iaSs1O
/sTmkSTCQYIyl4uXVuZ95DZCakPfkVT1oKtgq0FaMcyMmMNW1Q2Tw7odeQd3JhB9Q3OM9srWxeZj
vBN+WALmqCBo2dBc/e1hH6Ow1XzpIEPuRERAGTgeVlX/lrXHiZMRvvkBfzXVeaEeG4UD4yTJZ080
qLUYKWwJLOqthxKufj+n5IWg9o0Y9hO6yMt50sbIE7ZC8WyCXDTS09v49A/V1Dhk16eP/hFcwfRY
gdmCMUyAr6NH+NTyZbkRHxsg3pZI3aDyiIX8A4kuc4dehHh/qzIjVx4koraCbIZP7pLHr/U7XLPI
A6KWXU6lBV4oNYQU3EM2z5iVkgPNcwqghiMnRArucJ2hqh0AHYU3nmHY0Rmt7Abe8nUbPUSHAEIZ
Hb1TA7mOK5eIMNEKpViwvGssPDP1USYDFjcYDVunx/8M8Sm9466Ub2l6hXYwUtdHQ3CIaehStoNz
JxHcHTcJTxfpB4Mc35mqLKHGoFGColO1HaiXYbvuCwEnHuJDM7Tj+ULUAW9SiaNpZPaLydS5ljQX
Unr6JtLAFeYND3YX02azfeYG84OuI5pgo0P627xXQXnJnA6VxS+g/gI1vIVjxPY59nzng/AmckPG
ILxloa7hRSwQBxmH0njRDL0eiCd5O8e42OkWpbI9E+KtE4dN9pODUoeGcwPBPCpNF3GRBq101Rxs
9uYQVlDcDwWSEsKpD/CyMfSJ8VKkUzEev79Hb7yD9IRHaP6SQGAUeOXcKsxziD7ywy6XSkkN2LRK
2Whdpx7d1s55C3zKGIRQmLswYNbZdi0JcLoBrhlr8ZoGb3DXYLXyGjIDKgo3hiMlqUmA1deUJWyF
80KKrwr9PisqUoiQrU01inYvjE0ltANQBQBhj7eNoCCm5VwV3akoLbRctW5TDwXZhPOYcSe9slIE
UwEJyB6/RUlH5q1Ui+iXdrksq9q7/OMWRa+TyN8D0WcUJjWMnOmRJ22f74RZDrjCixvi1uK3YBBk
vD/pg004YCiY2yjoyxpdeMfuncDXOzZSKQdGmO5wdTTDRLxi5KPG1alx/mYREcPdopFZPEoBNuPe
fGf4MivD2j+80+yRq4B098vCm7x2aRYI3bevohX2YYoTjJwUmJCOHS9ovubidfnz9ccx4RCUEjON
a5+2UmdcLugC5iJXpn4Dq9ZOxGdj7JVcltOim1D2aPT22sMWrDyE6j5Nj9RpBXYNysityjd3RgRU
3hrNBsRPZsinPl5KH3Kw8c3miZWz0c6MN5NtSY7T0yczI0iZwtbC0N2zTbSZ4izrxuj+6HjIg4hs
KOW0hUOLv7p5JosQdd82cO6zabkwwNlJr2GE5/w2szacNLfi1xpvj+c3Oe/hscK4SFnEH4wOwFxc
pSlG2+q84occKvELibpkDWE/7moc3JRa7EEe7uhdPyA2EPFEkiX7PpNzO82DzVgqS7cL2cTImrJL
MFuFrm5r3ID5xw0LRmex3z6Hkey+UdFXq6XXz+sF/ESLXuSQI8j2DCNNOMXzbggsaDCfOK8CTMpw
AoNliF/5ZmI+HT71XTAK5volQ3UoxqjtYBdrf7g0d/bmzbtJ2VqiaEnPCxMhLZV+qXwMkjfg1BMf
y1xc6Ol/OJxoXrNjzZR9FSl/TV38SxhMmBpL3olK9ZQy80jRyUr65QK5Ld25elHijizIX60DX/TF
K6IXcbg0svjU1/G7sudmtYPS2mo/5LRX97NG96VCdCJvWSjdHGeQ5VZA6el/ckohwK2bFZV/cp4w
Jhf9G5eYhH4yTQagUXzmV9jlTyBYNogrtGPCww4v0QmFv7quOGDEoV7fhl9Pq0DQM1gOt5/VWkdB
2ahiognI89Bqb2CHIfgkHeN6xR116wfoGIIYlQq1mrmqbGpr2TUX05pz7HDL4OkaxXTuCx4glQm5
hYF5ZsCe4vfw8plZGPttDP/wwynaNUBFtaaFQDt310YdbFLpwTzfGvqJkiMK9ifhTBhNT6B+Ehko
6dEUFunyI7jwywk9Pea9rVArWeEdAnZyzBZN9iKcU71Lmv7/YBmtFHPCFdSc1XlMXfhS7bR06rSA
e8dmTyLq/dUT77R/k2fSLgohudOpUDCrefAoqHLpwek92P7IEkPIZA6HOGGOm7SY6BooOk5JShBF
zGkink5+8P5FfFSZ5Am3UilbPbPG59W7DKFp+htlf9TNrEeZJptje/t0LYDf0U1BBLfXtc8W/t+g
a8Bb9Q56aHS7aoUFPSofdBWTK2oWsI6+G60b7S0hVFEWV2HbqFzqJOOXzlqy0/cYNnsjC3OGgpdM
B3/KOXnUxb2F/0peNRUBedIDwVCf2wYidkNcjOGO4WjkZaldS0lRsRvuVxcVHiBdG0S/KVDUmduZ
6AZBV3lyAJGVtBdAZ8maA1y+zntsNWA+FuYJF4fpPJz3fuEMQb/wAPuZ+vBKk3Xb5XG/OXt0zmYE
RZ8sAQrMG3OG9yxMVCMRTbqnY2THa4Oj3Ov3fr/UpMVbGPmhacmfpTSZcfThDvZXTTZRX2uBL25F
XY7125GzQQ4/J6rPnH+m09w6MR0ckmv54eNq3dE7YRjdQmu84zME/Ye3mxSVF4TQOuAL7bmVhmhD
aj5FugUa/YWzgujLSziDIzKgdeCab9bVPOFa+ndFXjGTzbscrLiquEikAlj1HxwMlg0EP+7XH9gR
sIXnSiNReZQZRReHo+Q6Sh9Zhn5CkgDrlanhYKqj4kXl7ny/Wlo5ftH32Q6CqKVkhFAjHBbovcjO
7XIGs5qq+QNVm91pJn/FG+fx6q4g9X5cdL4XNQtAedNPiz5dXJfXd6kN+rsvnrSjxnjSnBAuWXlz
wzAwyXCTpAnwUKPQ8nAgfCId+uuFdez+blNXJtFs0ZJ8M85xQvewA23CriunIWYqTvcG6uQMFggG
8OFwoddMRrNsPsyALTl/459S8MNo0uqv1SlzOh1Gia5YkOGkjMLAFa0tK9mAkvzFSk763l82XQ+j
oQoK5THGJZbGS1LO2kIlc7eLEO0Sx+tE7wbj/Iat8pkQF45uLPTXelE8DpWWqkRsYS/Z3rJytWzo
SgwVVbkZ60e46s+EHhI/b5wmx8+8FxEnkRU6qMqbmMNWaSh0CX40HFleKK4suDzb2/i+xHoTonqH
Sjumwc+gREW4GJrLTGoheV7A2WPvncVNChY2afQazLlGdpuiIfCXzW10JUkTEvQ9Xc1RTRmccV3R
H8JPBtb25hK3tZrMIIO5xmHpLrdR4FR3saMjyxcn2chSqQVVVjQ5mV0xzEzc15lzgvBa8ZV1po6E
PFCQzKjX5/sylWMx6Wm4ZF9a0U5zjDID+V+oFpiEcasbYaiP5g+3VvUl/J0RPccpPxfiKcedrwNV
2uYnlpZVkpTkiGjukNx7Ka2Wa3+x0k0GjkVskuS+t/K06jKlWkUwEzcl5BD1tkqtVPJR9uKnOqM7
EQyfcMvat6iRfuZSXrvluISYoOH8EkCkIO48/qlHjZ0/iPn2qh7LzlpwGCH+zpPFSKHKtuXm0uyQ
txKuAw/iJbr65OfWvSJKq6cdOM3FLXqD2y0mlwtBYuQnTYnpS2xZjWst/Jn7L7sEddMCT/UfferP
2cO3OicapolKutd6RJWSge8dl3XrKSbrRWO79wDT4uJ2ZIk2XoSgyR+e/J4YbR9SChniU25ujS4z
/bk/v5LvF10dYsEOzN0N9AFPnT70IBjGB1mVg4PXqn4PbBRW6E4dakFXPiF6Vm43mokr40Ty7wkL
LnaEmkJog6mmCCad8ODPSa7z1T8Sw5MPO6qLqoZcY1Xso7ng1NUqxBrjB3kj8+rCjkD0s1Apjg/O
T06vpQp/UzlL7gCkdGxTmxVaeFlx8+ijYVdJU/iV7A+XpvMRO559c8YhVRN/cVcsSb6tCcDr1Ais
gpFxFpYIgC4KvvnZthaXS7ffbqdm8wmqsyHDpX5f0Rh749fljnzwiuQobepq+0T6LhLHgW2BW4+6
Po6IxgyxEpQYEPQuNRdNcqZjkCf6kPhPp/xyr7Dd00sugFVIiOm57ljP3pRRAYAuuOCY504GrrJV
feS1nLvogyMIrlEkX7AqCWLHiKgVadF455TxS0V0U2e829uOAxL9iJWbuAfbWrZDuCGB1BseA5Ea
TMzSO0kB8KUQd8vO0Kpqs0Q9VbwkSdeXK1f61oDkt8oplydF0pDrdBeSaLDzRf6ow0BZkvQTAqTe
7ctxW8K+OAVGlJnM+Tsd0dVM3zOxTq30FVN5nCSxzV6CSKdLNLK3YSq2oTBbi/Iu2BRs9N4uY7qG
I3fOZnrt15btFhqkp+cwe9WiaG87tC6fAY2VNi6p6d5KBbPFq2YMP7ag9gSo4PeM//bR8lxFeLgm
6bclXbc6AaSV3KT+4G5DvKakdB4YN94QycHVHPrpGiHoxIFozJnvbLcL4Numwriq+NnT2SnH3bqD
2G2r67FbuabeDgGWqvHalWJdKNVsg6OvfpJqTJMHSk1tpEgAL3Nv+QvaBGKPXTNZvkQCV/RtOuHW
FWWwh0hgqLqTOZ56DPdaRVGDeZZajejI0aM8muBQ2siT3AgtJaWabtWcSoOgbrl+K0aNYv9KiaBw
eULHmOFSCT/MuG3Lsjs7lp+1Kzd/D53WHMpU3kv1m1bPZdXFevxMsEygnQ8m0jyQFFVjDCJKU20x
oZ1aLFD2P8nGYsUHpMjqL4W8xyyN1M0TTCaMSIRBOYxHu7cJizk3WZTFkpqn5IbeDEYoJ3UDtQ+u
79Z00l858BwA+l2gwcWKf3XlgwPSQ4l/ZNVU1uDCVwbrNN/TxiEpVA0ARIa1WrGBWx0nANjTjDzO
SMpyYp98MmGqqrJv9/jZMmx3o+bYUMc4vumr6MHq9kJjI612bOuV0Zwh9p2ToHaT6kQo0BXnjXNX
KYUUS/J25MDQhOLvgk0JQL0O8tLRW+Ui9EORPqr3mpQhLNrS6azYnCbQUG8TwMxUzX+SmRbHgxsw
qa8BEWhuKNZQtiKsTt+6UAfTeC6bJ2Rf3ZMIkoGyVo5hb8g8p4EOonZVhHfa874cVamX097b/qcf
dsZ270hc/tUaDXdbbpPaG4xq9Vy+woDi9uboI2nqr8AN48ycblTieVm5LKUB/coKRzRDdlCQ+kJi
Qfas46XTZ1r+AVYGaSPa0mDuVcRZk0eKimomeb4cBwBnK9V2brh/wkgoYYCQ178rfxjN9jLF/9z1
CHzFUjOM14JgtcW+XVd5XneMwDHDlI7HNOym/AU9QZUzIe07D4TGWiz0l9JhXMytOFAne2RQFLqg
//2LQ7DubrdUDXBhMqgB8rzpKjP/Z/nd25RST2WE1DJLMTxbFUODhFo2UdPH57RZ9apIxpGjPFpY
D9Disypt7SLgnOr5oI9WMdZRVNlU7PS2Qdrpk1y+Sl8iUH78osjibE8yAxaytiKVRefljE5Qf4EG
RkfG5t2q7f8HP2NxjzyA/y67yhje2tuYcl9eQWnuWCrJS8IzS0Y4Z1r8W1tWkicPCmfpQJoeGb15
kNjxY7IRrhu+OpVrIv8Hx6mua5rqbPnVpTPm0MttNl/fqiWOxCUYT/pVjnH2R617IXlVkv9hlV7P
BnREsJti1RIyQm15WqAVK/VYJUqiZBNuH2uw261Qct5OHbEPLxP4ETj7Rl0GPje2y34P1Y+Cg4w7
T/PrF65RRojuR21Xkoyqn/erIxxnSWB02xglvFTZyT41TlEnexwU5rZ/fS9lKCtonOoP0YxgTc+a
ykkf0LYVGHzsrcEf0z+74M4MWgCtM8dCoJ+S8yHXi4bu8EKua3CrfVTJHB3qW19RPc8DgTdsFEme
gBY5+0qEU6HTzbNHDPtyyR5p/KB/okNj4eQJweWHq7GCJsvyns+dPU5/b2bo2QX5dSGZF6v2rXQE
NfZ0KRkZ9Ga4MRRAtU8QUnRbeoWU9Hd3gDJBL6t7kKJjVpTPVxLcEBbIe36G6jYVfrF3h9TATtOJ
q5/kc90+WgHqnEEoIvGWEIS1iUzaX8GuOEKvbsox1tMK3oKwi/WVhbusFNIGNmZ9jxqs3jfCfMK1
8gWmR8nWXpeOUOlBQEuC6hOpF+SexvyMoYdCUz1rIHRLnUr5PDxM1/aROgtCjfNKcyRMR5N7UmnV
FNmAsBZ5OTVb0lzTjctnyT3faOLE1fYaBwPI/y8Faefej2HA+jyGtai/3w8fxRMKUAlz8ZcsGYmw
jpWAGM/dJCkL8k0/md1LUthBiw56bUqeoQ8Jk15F/hbHrPEZ+5XNF9t/g8V8ys6eXBUeRQG0PzNQ
3nFtr5yAADoO/5baFMtJ6lcpG9Cp1OdHjIHX9/yFoNdqz+wCn/4LsFfalybpSGEQq8Ji2WUfvWRY
yjHSs8qbRirLOUhDjSYNO6I51Del9kcbZJKRNsx7R+liFcK2FXYSPXWKyz7vAospoKeO5lnVGflw
yMGkkd61VELW2hcjr0wpE2O45HyvjmWePbDb1n2yTkdDXwy4+DGXSFcWiGY86JJvwKLGz92b5wpl
Ibt4mVgE7Lm/CeCdcP2hkGjF74bzfVG+eUU4MIvdR8MDQrb6twVtaHzIP0NBU9rO5Ua7D4Xarcan
cwOZ6/Pr7xsZ2utBNFgI67257mTiaP/fDHMkMS53OWniJ4Aj/SUnJ0aSNBVNmNxAwhcKfI+Uh9kQ
rcpvwRI3s09F1g8ohHSVyNeuraov8nv3CHnXKNxuvS2pMFbavW/7/ZKB/MmRkEs5LnShtBziyPdt
fi1K38GXd8iXL1lr3/bBqByZbqdwUpUFD4RlQ4uopdkDbaJ81H9TQMJ1llqmitM7mBSy0RXJUM6q
eMbZ1QfSkAtVdhcjXWvwBBGh3SZ9ltM5k5rYQ5bks+RRC56uROdh0WEJ+kmnWUdejmlqwAaMMnzq
m5gDD3neBejlCsoB+L+/EetT7M8Mj67pku8wa0o6y6w15skU1j3GMW6uME4++d2J7pES8wz/Q99q
0cctEAKAfXrFQcHugSfaa/7iKxqfZmsghTjFmTrUnRyNYxIaL078FLBcNYCjw/KlQ5Qhm+8qlF7f
n71e9+iW9RZVqnvz342hiAv7rBRnOL0QurU+28qgTb4FJT4NJZLiAvOoWmkVp7zefliEsuzEUyzN
BLZxim+qbQVQ55g0ELJ7Jow1OZfBdLhFAmZSgaiBBeASIbNLe/IUR7lkRxrMgM26ibRDki5CkItb
nhzXqhPNFUbLmjL7eOltevzJ2MTXFGnzsfOUXRKWp25CXh2cWyz7rQNZkFVGDw6BoTz222mrP3tJ
Yos4sD3D60BBap31Np6nMptf0pCipHzjGwIKhI2wEY4EgfI4l404Ou+4FULgkYhwy2jgg8btQcIw
NeRal1rtFX3N03ra3sbCO9jMoqi2fdUlV9+LIbQt60qmYRnANujTdb5akGoK8y1kuBnRVmAgdSqw
f9aLiAqCTMczEy+drDxxtnckQL1HERbpbrn/cHwuQW2AvbfymZ7odQ7pHrlAYq3pFSIAskDv8BjX
23hWDAnXRA9zdU2Xpgh+D1pA/rJXJiGdRRIaB+7DH00uX/2a8WQqElaOAj3QP1/pU6ZjtMmycExD
mgpRqtfrBF6O1dZYoEULDw03z5JDuHCibX92tFxSLUe3ltX4bgIZZnMrXSE3HHUGantdovL8KgUi
K7brT4sD7HEtyzwYp1FJYpgaJzKFesE69Qk6Ro/BV+tWy3fq45Y9Ht02u98876SkyXqTv+r2myqh
GYElM3gCXefXOn5eRYxyGBfLS1LlttAUog6YkHUNc3LrAvSsrbktFSda2/M9AjWCuWdzcq/RIBIG
eoMoYefdtITB00aPafAthnkzDdwPRfKFcEkTVRugUIxG03cvxKCMatrQbS0wfxko+gLW+PqdVPFJ
DwhDxopIYqRWuXp2tZ7yOwL8rkeZikYvQ5TP71bkT7+OOGlVKNUAE1guBtqiEHrDz89Aa563ycJ/
v7YqzdoiDTnPU7iAgrn9ezfDVYTlx6eQUKVcNBZd8D9J6Ac8wvHEouXtuJux12NmhTIuiV1m2y1M
1PMCMAshI4o7a6UNaGYrMSRVfu4USei2S6bMzC7Gcrb2Ol/grK6Y4gZKIoKA7IhPQDWaEG/LnCWg
xEMBTS//pIV7AB4+WLYR+JkC7r4FRXDN16toaPuJpVgxKI+gX7hGwGzXfjJdn+5ylmn1l+JXTwKm
BxcRBCkKXGwmlGQgmn7c12HyQ3Wns7sSwyGMzc7qTzIvehFNPycGsNpBSjahGd2vJYiqy5ok6Gzn
gLMuyJvBf1EUncsIy5upE2AUy05e3s5nH9uhd6WQhVZqQkUSRt7ktWQ3unNUNgtvS62sWQXE51QL
u+1eO6IT1o0YD1bdxiIT6WulBXGSCgN/UFCNYoo0J5XuM6e1tJyazfkB59xCmmrbWhvnclk8fmq7
NwEujd3f0pXBE1yE7BpViUj+d2cjGbNYApurYIGL9wzIoqTzsMlZHzoFgHlFrzn5+/bdQWfXbkEi
OeYbhkRlT/VloJzfZ2Vc48dtAmmwwDkQiiY9UkZD5EpuLyw2+kWdOqimdS0CB+vqQVIsBcEE7GQJ
22FwJB9P+M5ZtUGILV271zC8tkGlZkaZ5wE5s6nOZW79qwQaqxmVU59RvHXQanuwIMUT1LXG6Vuv
OBqf1qeOf4znC9avoJwRksKgijwZny9ZD/oNkUNtXIf6votUm7J1OAjOOY57FHNlj/gZPtIBL/Bl
pzc8TrkPOOsYeuKykpZCuDf3kw2n6QaiwiXodW4TtaLwShNHb5CsuN0RN4GFVtOHDjPTQdAILzpn
hsgXK4RV86KollViMet4p/ycObJqQD5Vb8AIhYCXMVMHk/IhT6nXrNGnqAYaosX7NxYkibmZyJzr
ZLP1sQxehQVDUeQRSXRewcQR6I7hZeHiCZjVeberfLJ8Ef/B/Nf3qlVFYfVjUQb2po/DKrZV48zJ
nJNW4ujQ9Kbe1EH2uZw8UQWryjZO/NB4un9PAlwljG6zL57hnAYW8Rd30mSLr1kBNctKndI2m9jv
BcOzknRE3br2edQIdTm3/UBd6iHiVhID3FOtfCDz2zYGb9teroyNi3RIZeoBVADsPjZPS/mdCHIn
tsPkdu73XQsihPrKKHtf7ea3bxnDC4LkNbd2CAyx68JE6xuZZljm6Qe7cJ8sI4bY2izK0Bzv7TU0
s54U93MMdC9Gw8CWvVHuKYOOkud+lzyORgYJxmvAfUgft8Edy2akHKg8Dph0VBlKfxKBRWMharzJ
Xl+fSdiZ/KMsIDlyX1dq8euhpo786u6z/xN9lP61zJ1JJuYcbBJ9L2ZrZa0ekIRL4xNGZJgOtSA7
vBBulv1hUW1cHJGsjN1Jmvrm1V+iSsPzWI6RU1eSGUe9MzwNikNbO0zKD9RDW+JfXg8mfnmWFKDR
VQ7QBMCzDJEJ3ePd6xhSaUAabltSK67zdnoZhj9dtIq7iX97oSLKGN5RNAvK7O9AgP7JKLX1jp7x
g5bwTD6eqlkVyAHOBYBcw1jqDR3N08XhdZnFOQNU5H5XBFlTnpe3qnpPNAE9oFpP5SrAedEg6mBN
LrzPs+qeYus6njk5X5hT4Lab6TpTU0pSHTR/bWGkEa93Bjb/yQlEb9woIfOeKOdKRa/84e9XWVZM
qJ+n81bXwuPMmEL4B3qpJyezjnQKxO2TBZ7WoC0vP7qyKtErRhwUQyv2Kh8SEVo/bqXFUtyMvFkv
NgsiggxD/ggzTY2NtCIhZ3vgLZGPg6Kpm8jlcEfn7/8QS2h2MC8uO9Mzn9Yp2F7wAjiKNNYW7/HA
YL4A7mS3nK/hpB0t89P6pj68bfSWT/RtkqkC9178ZiWr2SSqReivGaRj6rD8AKXA+1WjNoNblNhX
hNksIH51HFQ3k4A6W+/K1PeHvBzHmPPN1nv/ycz2T9x+FNnMG4WFXhpsfgWAYThPw3y318oFnUA2
2MHPKDCRYkBwlHkoXVKBiun8WmSStyGxLjzuXtUbfTiBbTO27hwVIs5sC8ky1YIY2LItKxZix65P
+2i++O/Q/Tb3JbHMptHvbbB4g81wanQaj5UQMmvo7DGb8fQEYohCGy/3ssGUXpUdJXXAcJ6lgS+4
Slxc8feiqfu7AsJy+hvR+QlEV3HbVNhJVP0DHNiE2l1WL5wLSRzYiPzkFPQ21rt672YuSzH9xspO
Nf9chi6QD6ZijJ41PryEFBcogCbW8qpN819zjxKga7u2Nb1IJu/w0cYz2IhUX1rAqFBxTdgAvlbh
OaJr4JzeoK+PSCG0VeyNqqt922xyCKrqQ/GItD2mqd7IBlFNepLI90KOIZvjIulPlZkB7JqDgDZ+
MFdu6+t2Nkh0lJmKJq0djLL1OCe00cEajmqNkWeuzkjIJyrJekORsdgQ5SWW0474wRKAIzlBCpO+
5inv6L7zrEO1tyqi7F2JWpm3ezAMxPkCwLgL+5B/WcHhzFMLBvBZz9SrYOZgKc11yTrzuoJqs7FZ
vrf71nOzwG7uT7cpYzT2OUeiyg0I/NN5Yg56FbULTMm6lvpfO4ESOwxL9F4+nVAJuShrX4KucFXq
oJpqoaNuDJEa9vkvnal1imlorfl1VNIyP/9qzN8zjjzG342YhUJR1dkl7disham1LXvVfp/E9cpv
Oj76BWXAVXowwM/Bz+MuYONS4v6LIdyaUX/KSDbFjkDRMtow1LGmRun3mkpm7OnMgZU1YZ11XLyy
SDEVq5JJCcwzjtnALN65WJl/+aDhLJ689+0ktTqKgSnK2SHadfieYI/uD/j6pZY6Hm2/mNPLB/+N
i0jSnFWD4wgq1XkgKKnWIGjnRlcyYqv8fwwTHTau6mlhWpDn+XBgi2dxox8jwyubDavOpiZwO2FO
0hrag7LcCjjqokjVigic3rMZcSwNE+5gxnnZ5C8J+GZElsU22B+SJ+d2vIbgSHWpyY2kG9fMEzLD
fg5nJQaTnr2jisEThDu2fCJxIe/rvYiBt0QQjI2jmCafGfM6rmOup0kYX2xEu8MBHyV6w6xRks9Z
oMIQf9MJHCIRujw4V3layp/G22mLHxlLenQqEDcUn4Y6xV385afzlqH4ce1AWsi2fpzoXTPzTQDj
NXm4ldUq+FQiuzJn65glDABoLl9sB+Sf98hJd99prkgb3djKPHlCK65ICgtb/EfQSBiXGY/wMFOF
ZhwsGVKwhW0hiSjwrv/VD0cnzdrGDaU3heME/sYWwErzEXr7z4hbzFwTibLUfdLs3IuJk+AKi3Xd
OQtpsq/zlG4zAPcuStJTr7f7EAZ0M8nqNxqeOU7m+/It+9+qzuKmUXYcSdiUOdpO5XOkjojtaZG0
jDDC1jZvVZRZv6ptrLt2s9J9xfFZI0H9Jc09g8JWqipSSAOcnuJavRq6gHMbbDupzfg0hDeIxkyX
zKfu9FpxzW1u6AWHwFHr07Mn315oVQb8RNdn+mbLI1S57ZZb0CRSSLT/26ogqceaS5I3K+6m/Bfu
7ivkY4hdOgIzQxulTS7cQq8gE4VK19HY8c3xSjil1PyeeS3mPWkM7iTOBAw3tkTX7B72Ua7/LxFC
5EoXDfty/Z9O4nUs0Popiu7+yCTbx3O5hryHkvPI+GdXTFz3fyifcq4mRAjbfFjH/W3i9OwQ2zqK
0KgKhTUNuXC73clBRF4jbVjCZKCb5ABGlXYc9R0EvwcFiPQZO9eoBYkyfKjYrmMIRLvNbSZVPS2a
Wyg5rgjot+f81kQhMuNtbIjc5G2BFR8B1kpzk6gj3gLgZBJSo1prc8z7gaPfg+tA0d3K1SIZAkG1
/qxmmqktouJvsrNleebCHwe4Qjewvd3MqneNzeWV0Ml6PIWPYzmK6/RJW33n9RnMc2/+Zyh+F5g8
gMhn9b85rTWshzBK7v1vrN5xphgHQg5x9ZMqzqe6rHbUoHvjwOsTSfaAd6BTEy0nQExaFnYJo0mU
zTUgnESgsEWWciXGnu6PGqUWovCXwCnanF0X9oVWj0nEFHlhcSs+oM0rylGlzbENSGTkU2mhuAkB
318WTpHSz1NTTOnBsQ0vjCTXx6kOYMkBePKOTfsshAry7FgrBoxMrx7Doz+8PG7wezXNY9QDld2B
u7gqFRuD+zBshP3m0jP3TVoyOSkMOR0hT/diKhZrjk9MSj2DuGiP8MkDrYTstBnkUz2f5B9yOAHL
MuUgZLM3PQY0tbm7Wt5LDroCdaojT05vi2DU3gCmVNNop7B+B/i4mbAicBQnmoDI9r/lj0yWEAD3
HDVU6PWXWUG0wsZDS5Sv7qUUuMbXo6rS+B7FY1j+kFsUW5APT69MJAUrrsBuTOK0Wsu1l8F/LBTq
oB+BRjtsxhOHY6vX3NHWH2Mp1PHpiiw3zxQ1zVD3W5DSY9Sc8Fpl/6pDAC4J0FnrpaARrdnKlxvF
nuyfOZpi7qciLs1xGddaFwDD8AJXUG9FRpYDvNVCkfxCpC0dEIhZd1zS2gxS0ShtYMdYTklyr6zx
KM7QwVqlO9F/YatPZqaFx0+69uqDYhS2tJmyF/kdWSXHgL+CKO1gqCNc1aW9gYCUt0kbg6AOwTEG
56lm7wAtUn8y85zAombQq7lMu/x8ZgSaMvAScPFshaBhgdilEXaQB4Ik7b++vun6Ds3GoAJ4II6X
1Vng9BO7QgMYGwgdp7gc5eyt3sMt5tPO6OwtoumFnw4uMNhdmI5n/arjcbmOeizma6kxsOtqT8Gt
bD0q0nUhjeIeksfYUk3CZj2T6HmTez/TDeRZez+w3BR4N+xL2dkksOJ2D5BvPzhaL77AAyoSi7An
pYYIVg/FCV1tosKdrGqnwQrC3H9Pgm0ESmZgzKwi52vH1KDLXpYFUqqoFveXKyNl1VXk1ObC33QC
tHb45gxf+yZ+0YziUkJZZV54L5/B7XrSOC8DjhLJK1VkAelWsVFOi7cxp2MxXBPE2u8lRXMyfYN4
WNb+ldS1UXsGnPl5u8cwJT8deGzwCI9w+Fi7rFQoNENs+S33662U3z0BE+zzT3Z9HwRNyeDWj/9Q
AmPBvcpoh23pBMUm0UEUSwzKNy/uRhn/q2mhwKphzFyHGihwaI3itoUH+dRIdYS2f77X0SXuCALP
jqBsOVrrPvbLSGKJEwa2UVnfzO+eXc4jRJ+7nBMXL3RqKb/gBDT0oIk4zaI4cqGAHGQdDUXRKEoX
oyjWzy9juAhF06wj1urNeLltdBC6nOtlmxEx0JtJIlcDpxufDwGflIYSYnH2AeRc/EG75xRR2yKt
FSnQ3DH822IV4Vzwq865PbRpwGOOaBAFbLO09fgjuBlA3cTU2K0ErYFZOc2CIREvziyKpaaAVm4d
aEi1GyQWM1RvNzClnMrznsHN9pBjDvszwrnEpN1kLPumkrQA1S6JveEreySoReOcfDMq6vV1aVit
qAHCS3S3LwFRgfbgo/h5L7xs1yBISXWyAka23apIKVoSOQ28n8UW7Lefdyk988LwJHCohHT38LdQ
zqmcIwhHOh0fvC/N/8373OATA+lgUxovPIWxrwBAmP9hZ0ASeTN32M1YgBjLMhFWtMgc+eLsqwBt
MBaVwlqiFRml8LYDMESGzvitZf75NnpKMkbddfT92Y5Er3fVxJgaEdScEQw9VCUPd3NSEbhVqgCm
Jn3Zm8UeM7/2v8mxxAn2rTplbfhK6qett3v4ZjTXFKt85iXf3mc2lx5qgxKBcjlGOjwu4IJpH3gH
ULRIu9wGLovmgncLSVA5IB4cwU2jOfwP3YUbnUnh4jDidTYVHtVX/gQyeNwXXMkMMV5S4OFTBLGZ
aptTGFjO3uHmE7KrOOlFQPjFCO4Q0ea3bYhjHgl4dxtmFR2zuHIZ1yHOVPZu4LmHetMeSInhewk7
gD78T1cnHljeZEFDb2vH7jsoIJftp/UZlD2xRjr1YZhnDA4bHB5Ojuu7m0EYyiROnVPcGy+7SJcz
mTl4clvm/ryADuwAX1gPPw1Y41ApurHM+IA2NmUNADHgo9hBRAby4q7fpcfWNZqZwukR8FqPYUsw
KLCEYNZVCPa0kYu2y4xttV6tgV3xmoGTr4WbRIhNfG9LobRYDZ+XGa4cCIz6/wCTKf2RUUlAmRzD
feH4xQTDCfJkR1Kds+UiQcAaJZh1jk/Cl+gi+wGnlf1YJzxsGHbOsGLe4L9oEMJ7TtStbF6iArEB
5qOxCn9lsC7rdvo2pVQaGucI9QYCsusbnYRPmjgVben6Q05IgBab3EHjZonnhqV8+saTAtmVzoQy
egs9RBLbE362xkoG3DATkS9/i5YhFPgt29R2WosnskANPUU9fsYOemRJjY3Xjav7jMd7QDQdf7CG
PiayEtFFKGutL79gSofFXjSFviLSnz/efd5LTMu7G129vc+2AGcjS9LUI6G8CI4uMNgYd5amt+po
j1FN50TkVwxbjQ1ao5AI3BwaogHw0oxz+IMYGY+TF+ObIj74rWxMeTkhCbr9QqeaiLNNeT7JToor
MIGp6tWxVw6LOmzwUxnDyOA09+celcdoCP/DlrueRMs0cNjgvP7SNqGAPw8YzKeozy/zvqB1rKte
CxNOTMZzYxwaLIdOFLx3XaXXSDzkfj3Krf8MPLxtpseWMZtKE3v5PlElx/OWWZI3HvlbGxd57zzJ
OqDQ5uNCXq7kM8iggjOHBgXj+gK+zG+hKkGcXLL10pvrsC5mZZfDRu6c0xKlEhXX6JfiMQfpbxhg
6Qb/Cnsv10+pJpPCoB784LHdGTXRT8PDUwlF+/kJmaJEFEwfsK+dvuHwx/86aGwrHo1JGJxKSajO
AqYORo3o9Y+3GXf49EOZa41cgFaJjsK0heZ+iSzvOzPwCICRSntSO5QeBOCg4sV7VyfU4UN+9k90
cpbifp6HVWf89FfCUEdgAtC0O2l2xZhLfkHuVL+xRV5a/LaBJXCBlQGzuiJjvKm0L8ettS4bBVyb
MTTzwZwRnUPIYYCpAp5+O62Rxs/kcYSc9RUr1VY3FPTfBZPEbJbtYA2Fum6HOEeN7yLK0egfAmsh
4xP54LH55nUFrh3dmap9ydNVGV7vvgx0Kp4KY72/PLEoBsZ/06uHKjeF4bQ/TBQqXyiCwk6gGTKY
0EWaCzgVPJEF5HwKklb1mGh/aZAWfvMFBP54xnphznsmWiv18+0R7k2m7ThmixoRrirIjdPNarV0
kB/sZf0uCNBciRP/PssZIMyffcxEcqocghkBet1S2kwobiWUY3QhNqgzx+rPAjjmQQ4rpW6CRmZy
oS8OuYulIy8ZkivCIrQKY2cC/7ci1IF9Kb9t0GEz+vMJr3G59zF5aFxktMweRAtglryYytb7pEHe
4LPvSLMbYqYqduq20mRevKLN3vbsx55V/tTa06VjNfCvE/P/d3aFU+QkfWiFBtIcwpcdIfZ37tnY
gC97NZjDO3pZfhP9KI0BglRNpRMlWxhY6AFdEm8cutkzQpCEV+gg55EdV0Yoda9C4a4BZWq5OBsq
0vJ1XF0XpNs8E+kXzSsb1AaxdUdVDiTPfITQL395QMUdaUDBoI//OVnElrhbkL79S+7T/UNBDHto
+HtFENwkbZdPmti5QTwHdU0XE5Zeg4gcjPiz/4PaPoUXFfLhjo8jY8P+jfXq/6m8j1NM+D3tBgt5
uRwrTc14q6XKAaYzKvLw2bPWVwbn/RvqYAhvNq56swBrOHjgXldkKQWe7qDVDSoM4D8r66dWvN3C
HvkctRX/XgUL2Rt5xYp4D8KR3GV4BrVXFR0cvtNskojGbOnUAPE68DmzfXlgk0Jqny1dwSTI8XOv
XtGoR4QDOqcpB6R7eyjzIlIiOsp/KusvA4xNLSlqpRgHqj22JKfW4L+x+2k2Ug4EJ2OZEoqDyRNM
15Ei6BJCvW9VUa0RfThkk5Z50YqQ5EQqu5ib4DnT5Hy17OqnJOxM63V0w1s9Hx8M1OqrEXmKOEKk
0YFxtIajvjUe9LzzvdVcdRU05eJTQ5Ysy091s8QF8XaATa2RDq8+/y4mUuj4Zv8LraFy2HkQXT4y
2OVth4C0rI5VRqEY5ze/WP+Dt8hfhOz+omqoLNpAhnnO39xL8fx42xkzVRNFSsBRS3k+8OxnwoFL
dPjLX5pN7Pr2xsLhOhJyP64ll0HdmGvwAU3Y+2ORxBG5T+iJ5iwvgEFm54wE7dIPhTknN4kS9Zce
x4oY7iVd2NwZqCkkHjoX4h4GM5Vh0t575JBWed/0PfMn8INJR1mqQ8NIyijuugtsSTCcrXIH5esO
NSw9DDqZa8OzgS6qbntZar3ek+7djYMOnvmrbA7d3ydn0tcfi+KKCZ9Az74ntC/rpwLYHaQ6V3xW
Ozp5lZ5n0BsSoDsXG0BrDSHrBjz+j/FwlaAQlTJQxg1U1dtLiQWgwXLbd20ZRjOUXX1GjJ8t6YGU
oZizS2XsFJAzmte+BwqBmCLNJliCXYBB7OzlyiDFgK2crsUqtadATVKr2KIzhLMJVjy+5b50Re0y
cGBdspPFWHSxGHOvvG/FG2MkZrssXXfz2HTGoVrwf+4FswMBF0MCy5d4lA7Nno7uupzBmBHE0Pe7
G4k0Sfc3rDZezrW0Jy88LJ5aoLRW9On66dyRpHmpekKk8QbUb8jBciCI/c5AGVV5Uxo0A7oG8F7H
sKbkD6dE924Oirg/FVpnK/exlwoBTj2OcYUQGnFgStVLYkJu8S3bkaFcfPkDaBx1hjNcv6ds2ua0
4aQFad68v1VqRAprE2OlGXBykvkkBtHIjvYe4NCOSIvUJMu9WPy/Q8LO6/UgyT6WB1V81jIn5IxU
69whujwmcp75YfMwNhk3IpcYA+eDJ9Iod7c/zKltA1F6CTpNYGAYlmuz8JAJHEsk8QGZRe1bisne
/4/tHUyyCNA1mJKeyo4QiQqxRKA0JtKmxlSzecF0Dug/b4U15wjJRalnujVEESgBo9CvUavYXRci
Yrd+2/keGylykwE5j5eFgQSbD2c3WcPtHx0mERKQzrl/1Ydh8gHKY5JYIjYUpgzLkxqDCHcNPiDN
wKqs1rvB/lPYt+2k9QSUGJa4xEINAPSNFG+EPfdL/n8YjCCSpQZvp1MXLUAbTqoP3rRie+UUAx60
7jMpXKkrOF4n1MLBLsGhThxJm/rSx73H94f1ZtWci+G2EOqEf8XtrwVswk+1c10eCCo9fSv9SMGM
4gjJKr0qguECs7c+xovFccO0sfrNYKB9c/si1DpSIOWhVQeVndTU1knxqDov51lX24jH7fyQUCxE
h9hn1uvtgjjjYFHs3o3Tn6/gfbwagnAjufl1rxUxm9cfZQ3tiihcEWBEWT2LBLs583yLVwV0SV1w
xqKAUzcIZLPYdv0HbRqi7KrS9K21vf1+otvX72TcS05T41/2gNdyTR5FTfCunqSxvN8zVHc/Hgy/
/k9K2nGCk3GG5XSp1NEriROkURawE/t3rTMX2JkyK3d6aNE1uz9uCo0drzQ9/6nms1xE/47TzYyQ
5aU5K1UVR7hRP9OCOha8V53YR07ELWG33RiAosyFef298EwTLgeMRczQhXe/Wr4xhasvtzKMXITT
V2ZLr223x+2UPMR6LlY0Qj2nGIwk6apUccUC2MNXhPvAX1STzioujgpsCii/ITAAkjochPgvuZiU
fiMjz7lv27DZGIj5pVyCWQCkyL3sKGaBmQPxewLm5EiOTf9Ltuds4FLW09bwf6gQzsooBxb5968W
ibFUs5wjGxQI3h+HWDq7w7nY7QUiTB0XEQ3zk92obeY/8a76gOrAV8NoTcT9GyehN88x3HYHjyP3
8pNXQdkefXvHMX9GGGsjyY116o2SVKprw+0F84GNqE1qLbVNluNLwFnIzLXTiyedsIcnLmR0hmIX
Sar0mO07ljUPhl1GaCQBBnDAaBkZK47acPywoLfRBcbmRtgEwjnQ6fwQvv3KuFce4vKIyYon4/Sb
F/fXsr71GIq/TnF8nqEGyNunkkCgJmjPl3AojtXuuy3w+2KktWIzIaDg6g8uH/vnVx7DFxJCUVCA
C6Oi+Cz4BK5mSU0y2i+nKYQosmEQpv18A5bxPrW8R5eXt7xJAshei1wwCtIuBAoxYNLnxCtiBWBt
6uncUS0S+SMseuZRrRmi67cFfKVFTfFun7cySB+Eb9Xioh6YyAbxaOMSd/sUl9LQ8C6rB7gMu9/T
VmukIewtfJ0vl/KpwnmLHzi/p0gHUdYmG4YKZl0gVI3I/AoUaJJklB9LrE89JNHDxPrd0NrS2A66
ILDb8Pp4tXCQy6RNDO/lPX35FHmVllcd2yHA1gGDU3Ilc0PM7gO2Y5bu21LSPX3teTqsO40zFTgR
JcnF/5/sFkjdJ8HzXSdnCgeTEq0xtdGuezXm2+lXwo6v+a35CC129LPSwSICAhEvN8uU4lwVd/GN
vB6kEY0wP3lb37S+svT2Tby1Cj+xkDEkMPDk2mURJ4ekkGhkCRkBKDUD/oNNjT9QsriW3oOPQl3u
VxrSVi8rENzTscEJHurQqd9HXck3DCMz05vrXS4TJQMmc0KFFmG0n220cvcq+KHvd/AK2KddMSZI
aLIoZaFQPQUstujgXLYxSXqc4l7XXgyZkxYuC0uP4cHEdAomnovpGy8L1dGo/EVqi7FNKD/qHvnX
a5JyB8NKsCLY4LYzw2/z+DlNZQWiki1Lcq+eBTTN5zvaMET0TFZxBZOnkbrPRU9W7yzREOFd6Ula
kkPF1PBgriU364Li6i56VidRgE+A9JIaRrEjHjeovX3fqmmpPMJDTONCKdZoarOGCO1Z70UWwWP8
fh/W0r5lnFqvJb34fdaSFs6fBRWcH/MiydgNDBqEMmuaIDkoKClBNNa47szyHZn6dTSvXeJRAWjw
8sNiD8+yoKoWnmFQZcbJ5jveWHbM3XccMZJrvOiKj2L/mtd8DgBEViBPy+KVYGgZwMXWZ8LXxV0L
J1rP1wrPFsC3ayZUfQQ08NLgKzpFPoFiPyACPgP+gqKuRJqqfIShRhtlHfq+c4FV/xmEGkPU+sPC
RQPkWMd83c7mSyom2iBW11Ps71Jv5dtFy+imbxgN0+e274F1wl4YlLVCo8JDx97f7TP1fnp2zXke
J6ZpnFSi+jcwnMvfhtMDOsSvTVoFcBxgBrCm3g380A/BA5qG2rOPCReMyAONeV9yjRReWQ9V18tF
766woyiDJREmDx+j/gJAX7J1laWiWBYOi0rk9e4fgMMR4IxUa5AABvk0LZBBwUjhfN9Kgujn3Vyo
spXyoeJxjpa3CzeK++QRkR81CDKPCfgQL/p4Bh4q4TEtruxrEPnyX8BeI3zgX50HETYsHlSGOl5R
ngVza6HrpEdDvEMJclNPtuavxrHLqd4UDi09dE8wyfgv2Aj6LvXPyCfXOWQ9UrD5YssHzO2qyjyW
mYJAaUGEuMSOZ/i6t34uam61KGe8/UdcSAnc6fMSlbuNeH5Q469wz+sqawTXJkwczZJws82C+PPY
rVfP3WYWJEUW0flYx81smrs7lm74A9wY7iOjch9h8T7MyIB0wMb9W+M6/98ml9Yd1cmv3A4Z32do
Dcq0YEcJ0y9IghQrZK+IjAgMHfLl2hmCU9QW43ufTHPNBbB1H8QIj6nx3tK3MiDtkF1ppHHKcULr
iUkNRON6STDY0F2LbxLshXDVfrijeBAenOwUsVEp9FNhBZTLpuPxEPKkp0lUMKVl/dsR3SNrmxqm
VKXW4W3xRl8YTft13YEdMvSFhcOhcy7telaJJHc3sJpvq/JYU9HTM62MipjawtYb0IJi6gTFc9wu
bAtZJhAHCDVpPu0L35UK31EcXjYZ5vDfj1OdzxG4fWE4iD0TdxGawaeypsk5wefCPYOcpQv9OTWB
OWVKUJCWawWIjH8MdZGp2qr9O/hqcIN2sAYu9Kyoa1Sp7/GU27bGXK426t1n5b8Ibdrcrs0S1QQE
dAqbAOcfNHcJGfUbjcSoeQ5UNEkTPQ3iLVvptNB7INHT5SKqdKXX8Cmcc8N03gHssrKyoihfj2kq
lvFBchZsAEdjnjDUttE0C5e+v68aFzs/sCbUtLb6CUWFG2toUyxOWVTSxkKJtg+O0zY0a7vjOtBA
7cVzvUuyD7HitSG32rp56U/VyeBiVXRr2Er+td7LmvKx2+EcBypDoN04wdN9WLS0notopoypN66C
TAXFns6Xm2BRoWhSAFoFXQIdiyGIY1A2z+vToNauD/5m0nZMddlWY695V9Uf1Ri6K46eSb8DJ7u8
cLH7yh9Wm81uEQSRaqvTvtaUEGk2NlKcJZXZUh56BRTU9BxCSAkbMZNddzpwmqRqxK5g9dyERGkj
5dahrOJ4c2y93QucS0HQ/WrOOupqUV1VMwD4qK26lrBBPlDwGAopzClRiePJhU3nr+PabkZ9432/
J1WbTw/HmiUmcapFne3E7BOH81S/3lK7nEu28AJoZ+fE+mfg2yZt+4uqgSsKc5TAexm5GntXuFxX
QHew8Z1qp5dBVWIn6lBRB3VMrGDHm3QPSoTDHycVyDmoclkefLhUPZBAzfxZW9kgkBQ1hOyABZAJ
ZcX4TYlQp7VWWGmohTMpbi7r7HJ2151KeaK6TZSzGkbIyym7Lg24/J9LYjSCcnN7iT2+XXcXfLnB
YmLBB6GaFVJoXynU04A5eC1WtLlVBxhoV8f0UesyYXTTYtDHr+uznPgpUS1KXl56P3U2r/d7ED/N
5Bbpg8SVCAy2qcXO5/4xlCqu9UovTnBsLj+fzv+V0x/uS26fqlL35t7di7sEF+z8dLR1ohA1B8Sb
WIqE1OFDWXyD5ibZYz8swrNCc2CDW7O447+GfBSwKQkYB9DIUoIm9uND4hucYYPVN4DbvTJ98caU
GWK4fyZLlRU+tMKlvT/8DJw37BQMfiTn1n2Ksd+U+dfEWM//CIuCWDlgUhv1G/h33xr6ns6b90Nk
oNnSY4Jypz1fqKEc0K+gPSS0mbZCHVoC5tEZU6HzfZ6rjIuwVXItyainqY4ksPjo6uUQr082fc9L
BsdYXwHDQNU8rVUwaqvJmLyODJqpaS77KjTl+uA7hWJ64KYAoOJNWx3MILUfsI0rcUhPEm5l9tGQ
HsiWM6X4mHAqYGNYTL3A/vdNouUTFlEd+ViV788AfNndvvAVC5BOwSr6cA2B3lO12YFrCHEgcWvI
MDOnueAWgdF874Zpi7s1367rBt1AU6Hucdwov+APHQSMzr2jhmhh9svQQg1QGPjJNql5LC5jhqgj
ZYwslP27ucI01WxW1VMXqRjE4K1P6xTl9IlfqKFSLK6YgubPAsC6mjd4TnFZ0BecGbrif0tBZEXc
qBAe0QyAJaW35wG12C3jwdjh5oLD5gmj3X0xxGYobLhhiebszoI3wiUKoRxImImzTdYjVekqHbiA
aUMieM1XDRv1TYTpo6MCxH26KqPe2fIablb0zSTmrceLH3OekTKtvWil3YUg58QLpR/rQsESTtZ3
hi20v2Bl0dmDma3gVjY3JbccpjOGefrzq5QTP1n329JLztrgwtdw3dxqgXYRpQp5ZCn5EUYgolNX
2C4I9GKygS2kKcjmiC2FumCCpjcDIc5Whdm2bsKRyvRqfukIP/jvLwy9866X4c+U6gTgf806lUit
4JQ8HK+4URMj8AEWneEnTX5EsPHFcliRpPRakJc+SxucJO8zzC3s6abZA7KzI7vg/BCm6erKFrLs
g2MDeoDseiGvcN2byiQopXnmZ5tQi/0GPbcRZlHmhikYRMTjVFL0wFByGGpgt+3KkFfOCdjc0Uc2
gYOqXpviGxvQ23ndJ/Ks96J7Y6oB5ANnsG5ntFE7CWrvcYcnhJfVCxxLlpeugAc6Vb3YXi2OR0YP
tx+0sfpINGbzb3A8yIrQWZ9JMNPeaSZgCXyDdT4nwoVKDCfP4VLAAb0ehCYyIDEEVgyxG7Y/MkTo
L5Z3YcVKpXFut0Jnv2ACIqj8V9ZwtCeSSgkUIs0EdO5q57oJx4ucTAeFv0VMxjgfiWfEe2Xu5hj6
H1XH80X1d9bmw/3sZRiPLLcV5C5VLW7d4M9Ix4dYUo6bkydKcu2L5nSM1dtNrkvUDuv7rsmY42ug
3iIhmZ9P1BL7WLiZcKf3FLpUG/OmsCabUuXTNn7HXyMVUkl6bex03aUK+Kt2uNh2isZx8s51Eplh
wPSYSUluCmn/lerggc0GReuHq/Myt28bzxO00ZEgDVeeVG+bcE+BT4QiUB4ZTup8gljHUXtdAQbt
OGfoC3M9paoOhpp98ctBZp2Ph1Ir7k5EkNCIrvSfpeuKF5bm3wN0DQ27/rsJTrXPUVHZwxaH5Knr
WE0fqasUOibfVTdpZeuAqy+FGE0XBR1vmQi+k8IaA4GI5Kt7lG2j+7z6ZFXRBx+zJ0wQ2pONksGM
bI04M6lJRSIBHx3YtDpu2tVb4oWlGUlcWva9+LT/bwxfv2QccJEp+Fwlip+p3mnFMgHiMfN6ZB5j
3BA5dCar6RZxvLEdlgTegMMibXHTBZzyG+DvqR67pELgwMTQd4wkFjeaF93lWRMOevVPJ2a6dGiy
w5Bd54TIjT29crNLEdzX2orShvML6sy+RKy3scd+DH2lRRitG/B0RH6VUqPdAx2UuN55zEIfqHPQ
0BuYAYI6+6NigX6gSro6O7fteoZx9zcQ1rG5qAJBWSvcBTYe5WnadEJG/xzpBGS+yKRXVDqHRQ4g
Fz9vXgjJzoQNX7atpTgtGk0i15ZtZciehmsh138putl2xSw6FxTZIArcIF2Z+ZgECAREUeImbYB8
u/IHDM+MuRmNM1/SYn+/xeZcQdqBwBD/fHiznnSEommH/SHoAeAdL2fKn5qfX1A9xN+XIuB9EBgT
2npqJumGCZIkm5lcBdfipWAQj6amftoJmlOK4vftIQNiN20gUemBodL9U95CcxL7bXmnnC0uxhu6
3JuDGbpDayyy1tPkm0b9nRJesVxj2R4jlgOJijZ175lKZ08C+grFVhuQl0WAZBoHkZVLzJs7Q1GX
F6KuxEQwo5yxwG5tx0GNcLQ09qLs6G10v8iNHsvK3QosQD97GQcIL3YDpy+12t0SovVvmKB8veM9
y39zQzchw7hKdr3fyQMckUtI6thluj57xBjXnYc+Q/BvYgitj/I+g5uWqVk/HKQDZo+UNPgwvKP4
luV4a7XQERDVCFWIdKdgnYSVrv4nsDo5PX/h0nkM7yxlcXRlNhuk0ka1Cqn34dKCBEEUeKKBXFdX
3sfjectsyM/nRwYbP69rpc4KAvHp6SMvGm6BtSHa6E72D0XS3Z+kcnEm8OqW/HbjwwnWNE3nJMT9
D0ospeMChPFJdFfUUIYKegaeCo66dvyJBWOV/Vq11XHqGIY1tN6maqvsrdbi1sqUW6Hg1ZsLtPN7
Jp6YI+d3v6pl6lzHJYi1ob7n2QbVZGy7RqtPZ+CELNIFsRGq95rMlYfErDEAnRK+lXBBIyX8CIw7
2M0ET9ab34HlZOUZI155HZsjHKlZfYS6yNCs4kDWrJow/bYw+fZfxHvIn25tJgi4fLuY5vEyZgKU
OGH6tyrGx64ejFXzCWFgI2ipgsCIZwZoj4ESRoiPNJCG5eC9qm62gtl5PWidQZ6gPer1jRJfs6r8
G4Sm+g4n/yuzSLOeS9iRxwyDGT7I4l1VAhae+g1j49l01x93znN1Fn9qP95B2PeuwtewjM2CiXC8
4yRdA/zcFDQJiR1wK8Ryc/6xBMBoB7N2yp9/QzrNfS6FFrrvBGnpMhN1kKvzTL5510UZApthxA30
W4BnD3aup54HbIw8Bv295Xos0aPhYolWiFkXPB+NaiPGJ1Fe2vl0DqkeZitSDEKIel453RnZl3WN
kqLD18EP7l9pOARjRN/Tw+iMNwku6DfagoVov59UDfoZ22FopTNZr7U5tP8wqd8sU+Kokg8LmzRa
/B8RjI99IgHDZCvDHRB+l5k1gSlAGHfCOTwZjTZB/W4A6Uiky0tA3gw8kJrssWLuGlv+eVy1fNUP
l4J+kZLd4uAYpQWQNfk0nNUzyhO9CLw/djMdh70pxuUjVWplX8rdG5fcmWC8RciNaWwxfE10G83/
urD/1/6UdXPyY32kmF4eZsHd8359APg/EerUy2XNpg16vIKcuZHkO67/4+OJvQT04zj22fs//ay8
RCaEW5E4nYXPyOYd9JR1eTEa42+8YQFIx3gKpXy4AuBY0TDYILIpe8TfQGVYGdbAshJgsDq4gMCb
0nqAXdLzTstLSHyQjo8P0MwyZtBKmBNrFRPFwA++XjB2T+ev0XEEkk3j6PYgQYdxD5/8zf8lYxLr
4QF/0czgeI9pYAvBRYvvrT4QQVrJSaxkKvelNwsYAfSjskUmYki/ql4NmRjF4FS1CTnuNB+ORUZm
XmxjnzJnm58TOOORwBSQ/yHc5FI6UpPvX0xipYkelYfayRep4ZyWfEL8hgLjOAl1NzC0F3Qex3eW
lANB4cNtHLqEBiXICA1Y/gRFDriFZmc66HiLosOUsua7zu2FGwJlJW9HTaQwltR3+nV+EMsFaPMl
Kl1xCbpiVpn/WKV0FqFCMHcbnb9/l76txO2bNUA6xSS+bg5jh87gJR6D96bw/DJBgUwZe8tNl6sD
EUaSjZPFdJ2TpWOIeWqz9txD95oNzCJdbDVeDp9FDxxcmDCo3ZR+0kmCz7y1S91iBCFS4TR/O8+C
D0I91MPdsjYJtM/Z7ZkXMCGRg9AP2vWrpAVCDtS13EgNTni+fu4KzYcUs3Ovm4jon5GoKH0xlazs
F46S7B2MNneA1vg9+4YFj3w+lQZo2DfIOCzfa0+Q1iT0Tt10gn9wHSai0e644KaiOaDhfRenUAs2
9OH9eMKxHE7pvYE5AJxwJqERxdnO3MwCRZQ7WjUeAfhRlt9WMIvVHhEy1CN01Jo0ueTNl6wZxr2Y
OlrXYK6AgWTxQ0LqwHTwimAsZKBckLWVcZnfgVhFlhR2Do6+vfFLyQeKDGJ+qR85n4iP98JVlGLw
pDaW0Jq2/nm+P0hvE9OJ3gi8RkFiNM9js0wD24EsZfa6Wv15Si1pyWYeIKtjzWAwJS51iIL+pENS
hBr/3WohCug6vQi/DhzLlBFzIZWZOUU4UeYGB1KyeBoMVYJM2dnW5jZdn63/LOQhxI4uQSLXDXGA
p8tYFeIpHdvhhUT6ZlH/7LtcJq0SQaAeTxEDSCVvNEZPga0XbcPgiAXERb3lz6zNvI87y6ygJCgQ
U9VYfTo6fzR9nWqnuE1jcT0CJBPgQ0wPVqvv5/SCZeqiMLjTRVbwvU+W3wXX0C1XrIOnFHGvU5Xo
RZFK2TdKik29TTBTLhpsR8MYsks3jJMvmQ6+ELR2y7O4wAw9biWLxtmh5RXjyH0APBk9+1Wz8ARN
ITJfmuJr97MdwFdas0WDXytxs37hprdPnTCnd4lJxX05NC4u6l82nG3i1sKmAaysJEoljhTB1FiK
OiTXfLlCMwJNKnEiuR5MUFjMtx+IQVEeLVop7HWDnTb2zS0Y+yy52t3C59fEHfYK9XtokWCSdT0x
gAG5Gqa3L0MNkz1jnRpftAXELupqvqRdSxqZKdSaXjMDWCBlZkK8UercMbIZYUzYw/PslVFWfsGL
E9UdtwTgTGmhAItG04HDmJUukP36tn6sKXVLy2jTHOnVfNnsbGAVbEsCxvXbwqKIGigsSABRzPIm
EpnoeJmhp79AawVe7akccw/dtSH52AcZ4QOD20UAAu0F4Iyxh6USOJGlaS0e59JKJQm4oFPI5Zqo
YpC6m6BXnB79kp6nEHunxfuxs5SnDLaCw3ofwdqMKmNmHl+zHRBh3cPvhfdRU/1mofeFcA2Ci2Mp
aBhm+HvBcnTpDep3Hw0Sr7u+Neku0mJj/i3pnwsWvFHYNaiEiOdXW+cDpx4W6BVXFfqTN95bSQsm
AKATMW+vu78cYkVK0EJCeijZeuH0ey/0oV1+OlW9id3jqrD6J2SgQjlr1VVnJ+z15qCBwmYi6ULC
gfsBCfGvGjPFHFjgNqsGoDJ8SYrlPu2CgWjZEshPd1iHj5Gwp/24aPjJKkyjPQrdlROQHsdU8r12
1YuPPo2hdqGQD6g/byj6BazHv3VMcUEmQFQJmZeKQAF1kFsqQFdZXc0qpu9HTz6THBxLR5WJq2Ly
rfvEQtpQiYLiz1ucZ1veeeqn0GkZrRe1OvaPvmqSxnonDZpm7RvYoS+D4mDHPgCNZYvIT/gIx238
boo+gE1r/DjR+oTL05bG3eWJBBdDe3aiPk95y/DfPTHuIqM76Kc4Xh2Z+WYmsKUSfWoc1fi9LPGq
e2/iRR1CHWXVw8FbxX6DBanjmO4A7/Fqcn50wMH5/UpeROL1osIOLfgNhF/tqkOAkOLMycKDc1aU
qvf5sW3wVmSq5HtCHrTqJlEJeziQfGHFsuEW0v15yUra8JkcUnBA8F95Llh7qOHd1TgzIMHr7lLY
vMpLDFmz2KsnFbfwpIezRJSyG6rJYTD59srsTBGSxhPdJcVt1YK3P8VjO3/X+tjmylZo8+pLP7E4
oSerin6saz/q/cWlh/RIwD5+rm+TYenSst1g9cXCxRvxSPC7yeVLv1sI5SErpYDiTs/izeHA8yW6
mXECkDeRCJrpKFgWDjkSOwp/ZzQDvgssLzFhF/nvVu/1ga+/8MDanE0ADyR6i65OiavQWSixaAml
UI5beRYRsfOXP+pTz9SKGuu8sWmrUnBRM6H5Jh4kQIeVGED5vRB985vsNvnOc03wxGcAOoy8VkfQ
LV8QrRW5a1cbPWzFIB8a8MwKnISHxej5wF814aIHFBUK9zB1KtSkloxlNtea85PPbLjEBmkESUxl
pvpVap3sOFYBY1D64kUw1HmPuk0FcBoyTrowyYg+gsPQ3jOEKALstvjQSJkFMJUZjKWAW3uwJxxt
jloZ6J+OvHtFRcqTawF0kSWEUQMMH6+SVII9II0+D5z4amCek16dkR0F8hVlIIliFF3gERRok9Ft
QmS0iMj/QmXPBfq3Itvri1fdLyEngqrYqp4K0+BEAWBKpzORZdZQWzIUHXzEwioA+LlRleG36C6V
/gBGToq3WAdCT02NsIkHX9E6bxCkj9K3i+9i1copz2mhVMnhbpNN2KpVDVfHwtfVOzWb0zyVFrZV
SEUtNMBasCt57pKUrdalA5SZ+5OBOcW5ApFvIKyg8kpRpdLpYZLPt/uCF/deijUuq3amiTmblETo
PN89EDHZRWgq80Qm9oO1LxGu1lHh7xnB8udkD3RjxwtTVoqA48lJorJOkcJu97uy5Woiu4/JxFq0
FoDofOBLzp3rBUxxVlylOQoDbngSeb6r/B1jllcfiWTup6woE2RPLZK0WN0s3JLwW7JBrvFlwmlj
eDMi+hqicDWYNepqoJJBCYtKBGdeIZyd2YkfMHAOqAoAAPLVnMsarJlo5x+PG0ZBqW/BS6PHHVSO
QFApyUCi9ZH8X1uPu37sGy7uB+ku0d1Ais6KPJMAlWf8qQUsGtMbG0/zUcFlBtESyOkitKEl2EaY
HCJSP9xj/+oeN73WG0aReWvqPS31+9TnxrKqdfPLFAwTfA2r/6/tQ8dAs/bQhqXfKRK4N6D5bdEi
1jWyL8sgccMgxCcOllvrCxEgd7vY6m3N39I8RvvieaAEXanEhv8yjOtf6rt67AA1xwzI9rkQitoO
YHlgMZujd/1uBCttA5B1b+MG8G0M9xMSrzXGqa+kMJmpdicJIbV1q96trR4bg459FqS+r7hN5lBV
33gpBoss+gghl32Fpj3Rs1z2RGhyOhLanNW1/qfyeh1qHCdJQx+oDELD3NPZTuj5TDoR/5ULTK1B
kHCBG+BzXVsMhJ1TjtQa2mdz5o6dKWmBMOgg+kjaeVGSXazbj8kWUI6dVxi7B+5EVr4csX/0Ij6p
gWmyjuZgxGs8WsnUZEYUImc2nBoDzvN12099wXFqggP4hmXp2dgN1fjW15qlfv+gfGEdBftG5ZaZ
x3P6PJZ+Uy6/p/bfySCXF43Tg4/mPJL6pRc0R0OOo/ymaA6JoQSmC6W4J6lAkoy7ZNQcF8nKB+58
xoPgT3F2LYxrXY0fA+2nJHz2s3I0/byZtcn65gXk4dvTXnIZPDZ8mzUc9pPZJMNTvdW8/U7LrAO4
nKE2xWwtvp1k+Q8aEPSEcwvGIEnMp/LzjfplzRg8oQQxtp/3cVjhQbtx+FUUEt8qesmT+GvxT6sH
zEhsSghflM7p8ErnrlZD841WtwNJYQnVTQjqFYiIMLZ+26u36+Awfd76wXCbawfYAACpon6YXQZf
EFXZX742G9yrTAxdGkZ/vSHozO5mt1RUSCAmZghUfSeVjfNqjr7pvuI1yfyQ20lua4Cb0DapXoQU
hNVPW5kWK6+UUdxUIhU6gOJGfKd3QHW/RLaWAo6siOq1BM+/kgsqmstfGOtbfv6kIFQ07761mYdF
wMKKagCuYzoLIEWrez6XInwKJxsftMiS5IhOWkQhlYWNL7NYqw2lRBuBMIinRkC5B2nHwW7sU7ww
6ShjkeQrV4rEtsEtOlmGnodwBsVQB0hCdmZbdgc9vBMQxaN8OLQbBiygB9CO37svbdUjyED3b8AC
fl6xvIgEUbwkkCzCMdpiILLdOUl7tnB61UuuB9dsNWyZoJL4hd31A9iZIOgwnx7u9TNBL2sW0gOf
itvJ1CTS38GrBlopl6fScGsUdbh0+dLxc2WlHirEjGx50bB+qel4lAWJ1jBIFGN0Vu+lvpAPZBg8
Vo/C7vf7ZDz+ghZI62XkgrlY1/dokG+oSx6sSRPaAJu1EqSrbUIurU6V1vN6JxG7ggrnFsOfe5G1
MNBQ89PE8SdzwQZIO8bPRDp9tHNzdJASV2yXfOlHZLtGCeEYNLCEXBDYSQ8YISkjrF3p6/OGBKS3
UkDfFwgNBzirs6ruThrN6DLGkpTKwthShlBTXJ7hhSFxENVePm0CxzK//RclYMXKqGH9NS5u6MRL
AAR608mn1mEBLKQzvGX747mOrGrNjBMFjVTvxsLiJjkhVp9ZoaHDU1VsmYc9dNA4fjgPEx0GbPrT
Dlfk85ikCV1EWsEbWHKWKrBtNphVCaWWNxG2vGxEccJJTbdiNTd/l7sLTgEbMKzT6FWaIZfcCJKR
Kcc9v9xvdJOEbT3D3sbUfkYF9NFjKIkAYpTaj7TAbwzA5tokvN5et+qwrolm8iQYl+W2L8Hls2p0
s7c6x4SrqNFRsYbWSFrOD/MwULryFyhG/D4sIuPGIGhAJhBaPURVK2fHpxExd5Mj+AVVsRbgbZIu
ePSUZIPwsFmeiltQ5Xh1fQR1TpjcHo+C7I1VFzs6lr2PkaWHLeu3KzyQffzWGNMI1B43tOlx8bnI
62gdZRh2XZ8RrYeOlVebHqkpXl+muEjNyf5B1tg8f/qh12S9AFa8mjVG1Y22nz99XsjBmeAd9l30
SsXTAkMe0p+KP6ilftnEa//PTdo2z3cIJT/uLvqxokJX3tNotNCIjFqfEb0L1LDGg5FgOEaoM+Jf
yg0HGNpsKRDxZpABsUN4ItHB0guyJjND1Rz1fuTi/DMD+abK0Kak2wn5eSPgycaN16obGETYpk2c
577UlF+QwRv5JYEwoXR0xgSXQ8c2go1jaDHsUOv4PjE3JUhphYyzRb+wy7oZvUp8xBOC1780oie6
DFjhZ2SleoT6IrBcGirwarfrXDU+ks3cGDVu1k/TIYWD/Z2yOJuVsMqhyO+Jz+uBa/WIvGjsKL+B
YZUANq00GgoHIDkt5rnL2iPw8r+gbKNT+TUzgXFXiDSQ/qFwNjMbTJVcjZV2Pg/BRL9uiMP1AE3e
jLZ0afSrRZU7Tp98WWzTMYnV8ICPHjMK4ZwVLjlxwurwwx+Ej6j8W8PPjjV5HEeDDWT7oEvZbvc4
JQbQ682A5uhExby2uZ7z8p80rRVMlo5GbPQhOS/INtLU4s53+BdvjlsbvvyYM0wdPacIk34rYHwl
d5yoPBZQ65G5pWTq85ay7+dnbj/Kms3m0Ym3BMny9GGCH1jio/azL74VS7eEaYa0t3b8rmKi+KZB
EO2qVi+RY0vIvP5NjjxryNlhFfMHL4JKOAYHttIHUu3muWQosfStS/Jl5XD3NnONFl4WH8DsN3XC
St09dN+s+YnDTOTr1PRkobN1UH58X1mWWbsxAJ/p2FAK/kyZ3gBYIfOUoKqrREu6ws7TOctTQ0fd
cp058JPaWNUbayR5+4R3cuk79UmiReC4+vFxoyXdDjxSSRMIlnB3zMRs3SlskmiFn50nCgFNCGNx
7YiKZXQG623Fj8GzaLaXK2Xw+X7wEka49PHWMyELMVqJabi5UwUgolOdaBktKRxu+CVxVIsffd2U
XR+9sgisUnOfLFdnnHvV2icpQpEz5GougqMLg2HYMrGpA8yPgjg58HWNbQIGAUUGDBAF6Bm8ZD9B
fTNFwg1p79fkipKZ0UoP/7WKXG1NA5ST10YvJcO7jLAXLyvkkZWFty60I76dv/Z0rwGhU/KkZFMy
OVdAxHZd2LgFnSxLSZgstOn0QBsBdAF1UmTO5zV+/2twP+bYdjorZToTkNd/QyAh+MTx8reO+GcQ
v4cFH1gJQiK5zGPY9ok3DsQnD1vFtdazCyJLojEFtX2U1XtPJiEPABxZdp6t8N6N9a/cio6JaIXl
5uDewaux5y8UM+vwSO2ijKPx3r3M5JJ451Q25r1cCMxpZVUP/tIOO87jWNG9G6H5UyxueF8SeOj6
1lQjIMJQpkjRv7HO65Nl5a6mzl/yTSwWkgMOlCo9ffTkvAmpWsu1xTTR5woeSgoU3lJTcXR3kmqq
VwopX+GGtdRYJg2ni/lCwuQYuDggy19bdvFqF0ShgrAXfWhGmzJiEJbUQuz6vE55PQcDhAdLP0IO
NEZDzexSzH47Yiui4JFFX4Pda5eEqCAz7y8+vnPsg/T7JUtK6+Pt2CP/rfhRO4q/5LaSy7jmfjGB
Vaiz9x5N9sJaXAXs70stBkjRSQ8SMtaU79X921EQUiboDue/9NqRFVdreCxIXcsN+PSTjePQ7GVy
2vke06QWZo5h+uADF1tw0oBZkhB7Ni7+tFocaoGUskBgcKx9dLH8i/hsU8s4jfaLvUdflhJxf3lF
od8BnBgKWDBtPgJbH6hjatRoCuNUn4i52TPfSArLgxB499+fUaAmDYV2iXkYqJNdxckqEBwFiL6Y
fuksvlDUFP5+HRaG0AUabmNH1jEzArFFvRmfWOm9MRUbHkXRmvK0KYsNZn15S9SvTH+2M493zUhU
KLqF2xf6T8hKndu/AKCRUrL6ENJfFWtByzLRVR6bBbESSYyVcR0Ma5L2byEPmIrJNa8h2B3Z0ALH
b1wkaUxtr2BvRIXLAIabsHtrNHswjrs1QbPyhZnVMooxcHfsSlloi09CHWmv0SLyDOZ3yIX6yr+U
FrcDPw+Zt7zwt++mI/iu8xjhLUKgTcUvA7T9utXYnv0im4fnzF1WTrElcq/TWG6O5JNlHf+WSqdC
avSs5QHCz5k9gFnfKSH7ttlfiAwqjfWdq/J0wYlsSbHCyrl5z5vRb5xMB7UUuPIzuJKKuKYcxKgk
W9gtlYzVy4AZ4drX9gSZbb5Y6G0lDm9Y72Th95GkyQoyOGVcml+S6ehX4AZEFsJR6QyNUGe7MGgB
xCSXL0EuPy6P803N7RkLOyoZP+08/UktJAcKY7p+HOF5zIS3GaIKaVJKhwSySHF6hl5InNo6q5Fi
+T+VrvTBPiDQWfsCJpeTXjiYjwL/txXJBw6W1eBkg5w/9j0Leows6N6quQwaMfMPgCczF7w49Zge
KRYvgUP1RoJsurwByjruMq1/ScJjCYRMPaCa5TERyHfDpe0ezdpozTOCJy74PJfdTahG59jDIbNG
M+ktmiTAKh1VOWv7b2aX/vBbsy7oqlUASp1lRddY7OF7RM2jdQOIzLdvdDHUsG5kftaNzOQXLKNX
kNaWOlhQ3i65xRCam7EjIRzapesG03TSvv3Ps4qQZ/FBrNPYKVXm0OU8efEq3PgDBIwhi5/YAOwC
yRXYR29nxxrwhCeanGDbOsFyYplphK88Ggc5vp+VWUcr4gyAPxs3LIPna8zYE+hvtQZgdlOxqSiU
n18Kt0L1RVMXuFP0m9W0DMVf5u5HzXYeclqJT6tscCoKK7UKkcog9GU2E/sjmKOuW9kdc0mcDWKU
JTNBujnqqIF2mgk+0AwLmdxGtT4YE4K8Jety2QpbNEydSCtX0vCZ0bpr1xsRNcKlyEdXXlTS0eZK
bFJJ5qEEiqwz2DvYHyZOo03eN5+qymZVkLfYoVXItTdIPn3YmrlpxEUIZRIpSzWMGKJHRjkE1is6
Nwj0vqmdTpPRP7Hd1tNGzdJVVy9GVzs+6i/A8I7t25jdW0PFGS5d62kSPmmqZQr5EB8EaK325o5g
kNuZZoj48g6mKD8655+z4UII49fn/9NPPh8EQcD7ZLKNPFfQfjXUzf1nHeSPsNfRymt3eQl60Wji
m6ustXVf7lJz5fyShhQ3GErSm+uSsACdZq8J4dtjfBH01tUBxc0MlmWvXyV8pxxeA3OVcLXc5aSV
139auya6oY14zf7f/cBhwMLMGsUJUOoKLybKgiI9sFCSzHvOOZAuR7hFiZHV0vhrbaZUyugXrlWI
YBrP/Ryp6effnGKiXRcPWmaDaRP9I7ePywWH3szNlIZL2eKGz5CaooJC0T0oFnACczoz6dt75BGx
S87dmar/AJPHlsiMAi3p8ASoBJz21jmUjhKsuQWqwn+pm0A/QXsPY0dxc2glWs6ZC1QcVnSZmxiY
5Qd7p8Ku8v142OzfhdSh1BYpEmPBz4z0oo8YVObTEe9VdNZBHdU/76qie6aMF1Wg7on9+vBboJ4C
CqqqoJDiKPMGLaIVcfnUVW/DwpEwiaqIZDyz7/OL57Ags9cAuAKjTNy6AM/H+a84qCp6MrP4gboH
Q6byFTB7naWck6aHgvpjqaEZuOvyqmmh+/QE6hU1DnWlpxC1yHUL+mcGAYyLSV/yxrJTs7WZ8nIa
pC9IvOUEZGRZZpV+S9Ii5nay9FiQTiW5vQmg5Hv3ybw+dXWqz8DPKRdp9tyAI8L7Ybr/L1mur6ib
mcu19KMw7tGKd1KjZEqeA44O3+bPBUFeEXxOIJtyZ0lGVl9FmUP8ohyTAwVNpzw8YYoj8bkUEw/Q
m5UDZylawVmc+t3b9jeKJ6D4Y4oiuNjmvu2HKv/DJU7gHlUIyGDtwZ7HJqB5fTV5Sf3Inuc/6yRw
VCd1GdBHmg/WNdg1uTprQAYOjugEC7+wuK3gwH3ILqsfrva7IfQtNT4quDNidEWX2a/LFIftg9DR
AtMmKSUrAyMO0qg9s6uqF4MO+AcTIOXOexg+V5j2t+tUyV9ShzCJXYzq3Qs+bN8eIRP4LSRjYpMO
qu/85CKQs1Cpzlp9NVNJKO4BEi3yR0vX4XZKZPss73okDLuba1agR+5Hj+Lkl/q4ruO3JSuO8iqN
OKjqpZ2EvdfIHU9VoZDFCOL842+gzZGnDAz5fGOFPUjSxj8A3KTbP+GUOdLyB7EZ1Iq4A5/Jh6MQ
3TC63SXuIXlnvLcsqbjq0WPgQkVCDVUW/mrhq8+euO3C56j47JmfTzbbn7Qu115ylDMwJx3FDeZc
EenKZQKQus6LC1VH6+v8ub7N8EYT6fDscsH2Xve+XuodL4ir6BlSMVlLTeHxFPru8xCsR6Ekofsd
4G13PgQQCvG7XyrrQdh7gqeTZ0GjS7YcuAdXtklEoq96PbN4M33xvkeGtaewR9xQcwevZRv5G1ic
EfdKr/dhiZ8EynEtu1T7ZT+76iFpWPVcnuPHv4hEpvDbXAnfq3zevw0cvqMpIzg31E6e/QFqS2Dj
kI7PMD6Qcm7sPMwKXyWZX2yBcjqt4o+4jJYmZhYAOs2+DuhXn/5r00Ve5ma4TO3xjE6KGlqNsb6/
G0+b+DZtYYk5vo1/djJ4NMQVpFfb8YH+6K6N99OjKbf0/J4AgY7XevQEMI5iodR9FV+vMgjxdP6W
/RXynABsZtpnCThwC+GEXsxAHhbYptOt8EjPj5MMu8rFDseIDO6XcmeXPFGAl/rNG4d2KT0IvYo0
jPSDxKMa6g02M6RFhTtQGLJ+ZgHjW8OHUm/JIbNPThNaDdYY5XZ6PRQ3aWG7DmUG0JYgkQRQjuUZ
gdPumQwg7x2Yd1JxoVcE3bPhK/oY2rMhwBZuH44fyEp/02BqjgEpg8IKotn/z2s8ur5z6DzIrVaU
uaNzSK9RITcVO20D7ET1pCJOS5RJIeCIOebeOUWbvZz/nwpya8gM90Y61Us7SmbWtCFzVs8tJw4s
7DUE2GrYe5w5oXvz7U2VD2JGt9YOJ7jbJNFIbPlaWXmanT0XJZIrLy5nYY4NWas2sU5coHTJNpni
hsgKczhglFXhYXxzc1gla/LGcYrwcolNs5mKnjqf0e+yWPbhO2g+ZmwIAhgKAKY17P+yOwPFU6Lw
uAL3Zl2Wbtr/bRV89ZVDjNYhRJCiNvuTKRRz7RiAJG08UB7IdoSbKc7HfhTkBnJQ34O6Jg/oGEpk
iLIn9ei6sELiIuutQ6YEGIsH81yF3flXHqa+Gvf2pofv4x3h3GG01NwJmuncYarsXocHdwE3hLfJ
L3JxRngBkxpT8dNbeB/3kIxodkhCD0w9OGqVtW4Do1+zuBqJe1j777eHv4kweNHfdc4+WUAATl5R
HtYw0aX52kttVMT/hzU72i+0AmZrVyKJnyN4Y0GT39xcPPQD1eMCNRWv5BpEFhCS/p4dYMfIYd+T
cLJZd5CRi+AuhoijcsIEvTIzFdWtqbkCk8kUdXtBGqnAZEChw3kg+uZmdxM3JTbA5iAka6xZh6cJ
R7tQpMuk2HhMojwwKWT+Q1trCOjX6U2X5hMmpB+nZI39UkmZ5GB+wlPi6GroHpQIaY+6fb4/AU5C
aHsVOf5+1E3qp2HwCtm9BDU1fo4ZssMS2SXbL7uzKkwFHHtT7J8LKukTg6klUCOHWL+12dI8qKVm
n2ODeJwpHKLATAuHIkDqHISbM/qFgPXSygHKU2qQtEhf6xI+dkKAFUR+xgi2GQ5bhcR1NMXL6eKU
febVps5NeJuhyyp8T+baF5hZ/iw0tQd1RDI6e8JUa4LUUReiobZGkn2NzAR7jtq2mobQCTCmWtGC
JGARakDwbVoUw+LtCB4Cx8vvd1FFPQpcFz1R5eh286TyZIOYKKvkULaHW6ajGa5cIvuH3sn3PNOU
xh3VB1uYpiGlMGHhdHn1ADGqOij9QsuV/gGLLg2n4Eavk3jO046XXJFh8pmcV9fbNJBT5N97+5Bx
GpLuZZ3KsTwky4LVW9U2O6EpXX/7CMKxk5YeY84u6ruXFAcilHoBCPRQKU5WU6XBvNcrVb78lHFz
aYzENSq2GhIEa25QstAojR8x7mmdreWLY7B2iKcRS5A6UWTeGAvKWFOw+sEZhKyGqDXqeOypLcn+
i8ipTNTNb30k9fL9Rhao0mXDgAF2srgGAUDcBVWBSxZUyMr4RioabLOXmVx+PPZYFRwkwAdxT+eb
oYqiLMWHFc90AC9tURVxg2tb7/2v8qVJnPV84WApnPIkcA3qJhMIXppHTycJjwF+FN5tI6dPYAgR
TpHA5Ub1hi/V/hnueZUZd8zscPpKdIRKH0dLYmRBpx9RB7+blQD2U9MCaSxUdJRxTZvB73qDWCK2
WJ48OKhyD8R51LQgUMF16xYlD7bQtjhJCov+iU/BLK2DkgxU3lCt08KN2+q2ieexz/k9jVOAW4bx
un0hcYUUIDvBta5WsPsfro98mlmXkg/0kYTO1QmoorxqSWGiUzNHXzrsCnpSQkmCcLL2vACYRYJd
nTk2RZhbioTKDa6+1G+/cACc/x3geTCgvgV3IXO4sWtg3YINlsrJ5eAgwQcyOuuW40ANTtGS33Ex
1VJ30hHo13O1lGMssC8OR1/s6CyVH3A8K+WyPG6xfnuj145RMRwyL9XSvcljKZ9QBh8erzvOo9t7
+QqZxhq41SrMooMLHI85WJ9FHKuFL7CMcLKErNGNED5SMhSAQez18PIu+1nodqq8X3xmrXAAiKiX
L0Dq70DRrSEcDkqJIY7azznTHMY3+lrX7kyBXEjWzoG/1ovUxMOplLGnTsBJAdpZ4xBltf43Z04L
2TEKRtoz2yRkjHN+KvwBJ//Iwd2qtSqut2gKm38o8JmF7/d14Ojlv5J/guO8hHNoXu54Hvt/BGQ8
prvbbNzR1pyhU6hQG8yG2VIR2R7KujQSHrFHgi9YSaoKt1QSAIn4YJoWjp8pyEZ9jyTvNXyKCloo
u6LIGBK505UmjyqaY11irzsR9nYvjf8Km0ZAvKCD0KPJScpfVs/A4GDhAqFeXbOkchK2BGE3a3ZO
5o3YTOVTRhM9dT+kLPdGG/2fImUl8yJFyxP57NP8bbefYvzskEOr1oFvPCnfXPHaEo3Ph/pQb4d6
J/bwxRr5DwLK1WONtt5nNso/8bqZVGeAYhCAt8XMDUXuRZkFSGbI0IJ9dIGzvNeK9HvUYlmhQ8cs
s6uhQpNY2aSofD1ABSZJYLCeVtw+6QoW1sWk5MXLzbMy5CPB4M6AlFZtO8M5kZFzwyMfgpev0Pgt
7OAHADo4OCO7GE27Xx9Xt3wydKgrYlD5/AM2FDQxWC6U/s8TQEXzfTrA53m3zjs5T5L/AqJ+vNBh
oijK+LW+z0ZaWDz8DNNhCmVrcqfN9iLHD6ymwlke41m8L7Ju3uGjI4l1tCQT3CGHMHN+recDMnq2
wWLx/ORRuycd5C1pDDtoDozkwr95sIewu53ia9lRTAaezN6nxmTpqrK6KAD/fnLAt7in8FLsKjFN
bkP49VBZu4BbAiimEacLD3S0+wDZoVQMgrvWn7vDO5hMfLDLMNXtRcigGSpSvl2KKVhT1XJl88sn
hwffJuOR/XjrqAdGqjwieGO0crHEqoOQiE8m7SGCD5/rN60ErfG90MM/k6E2tFMhDsejZ+T2ycbi
MfAPcN39wyBcBo4Qp3VkChLtNvvbBKVU2SnmBzFhSB5++eJqv5TfgjaW6EE5Wbo4x3iFxcV7MalF
48ksqQgR3CgfSUFAY5hWIwwIGMcN2EzpA+5vkDmuZQdAc+cM9ZIfF9dDQnJ8ltX+9qYyh8VLrwiy
HVCrxLWeZY2falgr97TIm/pxgeJqDfgH4efPhr6epH9D7YVkMFBpPgkif/k2368w53Bjv7m6jY27
QXfpMrZOmVG2/SafatQ8SFxadeoU/SeIh/HvAaIhhKlgyUv4/sAFQ+vXqU8bwTAPKILDfTlcwPrU
VGbTyPCYBHkwTdaDCJtyDzE6e94LxHXP/JI/Zno53jdJG/zM02wyE/eOTOJHXupvtAY4zMYCP5EL
hAtIjlkweEerbYNWt8+4RlFFjcC84GAlJ6VPx7qZ37xTOJi3OJUy5nOEBDJke21/GuuCF14t7Rfz
NIpf3LgIVgVonOMYcm6rlaOvTGruDU6ddp/L3wx59GsF89E1VolNs0BUTowos/Mlpi7dqfXQr/xp
asch67nJWngn8Ei+flh9zyX9z+LuGJ0yAncXWV/aqAr8l57Y5dLpGdYim6BhEVJn+Kuwx7zVeQFb
hTo7CDRCCJjV4rHMywHG7f1171E1gosS4J32osrTR4dEZziJoQ5s+MFfs3rZjzqfChaVOF0HMquC
A5tDfLVXcxTtkzPgFxR5vzUITwUnt5Z9UWaQ/VV2mfXbeEhR+9RsF4EGIGLWZ4I4avbhVJDarVvI
mHA/ngbM0I3h2tz+Sfuwh6gMRFNX85UinIMTwrYf1xdgJQHaatAceW6IwIW+S44obhXKfVAlAqHv
eV19LyjuPHCAPoWrR+M4ISUPHZkGqit0lCVGkX7TuxICpTwlVlHt5eCfVxXgvQpZFXCsvC1sV2fF
PxrRkJmW9zdo6zLN1QVjYVVOV0VFenN1DjbglF47Ou9Uwyz6GqcGc3tEzi4c1XG4owlGzlWfgS1+
p2IHueatKWy6oNL8jy9BjhfRr0nFBPPUuDbuwFkqcIbgzGvdc09QJGQhxsOT0XVJ+KQDJrT+5u67
d4basfMMhSZ+wmCfsfcGLtOwjHfqGQjSAL9vXWZFH+lb79tb5vfF+F10rqZpNZhVZAzMQ3kiXdtk
32eNODFk9Bt/j1m83TN8KNNd28J7kfds1O3fAiF8lcdd0eF9hht+RHUv9B4gjOnpYa2iaDk2uh3t
XJoljvewKk129NBg3ZhpqLQxMxo6cmCqQGwrSYFxTm9BPlLeZ6j/XH/+WOB5Qf/7b9ZJAjXXstVa
sFOlFuoPH6ZtE1M98s57OPUUjXggHps7X78V+8Lnk5HGF0MIVvyL9lKIXnS+7gAHlX6CIrN0kmhE
26cZxgHUNWWISR8bOyv4oyL7dDdH0rQjPIuD/uAnEnQORqSRgvtmI1Rv4EF68RNicE270NGFF1qg
ayPj4ux6mgmYwYurR3kHv5jMrUpAWt3LCyKUSJg9K6sE0J8sKhC9W3EnDym4GJdObdQT6vu5icyY
IVZq5J3r92S8PJGAA92YEAfaKmUD25Q3GQOGItGPBOfmrMtdpi/14fX9nRQCjB1DuO7Y0evlDNWF
Or0ZE8Tf4nWKz1kLEAbruyaKrBK7ZajVC+0ODZgkfvsn133XRytZyFEPXLTh2RAejBuS90gES9oJ
ZDlS8EsDK+jZS23Oc6l/U2MFa0K01SOveCDeA1L1J1rHSbMD05lb5IE8UqYjSFsNj+hgUsqbgT9C
uBeAxtDNj6XObboiq2Cv5dbTRDvx4X8KifF33dbn/AlvpdY9hQ1qY4jeJCQeSzXvlMs+BC6GlXMF
McGVQRCBT9eZxHi2pJ/0l52xkcH1Rc8N89yUpVwoyUUsswibNCo6DbX66BQP8lyldA9hZWR47xY1
9+baqcMSWqlrAgJ96z8d9gbNrRa5Zi7ofXuepXjS8G2UejXPX06rsplJPy25AxSMw/uP+L4xqIoD
pUx43KIPyh3qNy0DSgL9I07oFmmrsdtalpTuaImfYwid1Hx1/g/Sw9Dz/pUpdR1j2GndacCbUypp
DNbsLq9pWp1jjJnR2RnlFP/SQVbS+57Izli1hlL5n+yHX6ol9ip0R2yt2GAZcXtpMSNy9PUAvxQ3
xW16sGQZbMT2udQp9tXYXsoPPuN4y+WB6jpOgRL4n20USIhZD/g02kvYkA/YueHKErTfIrNDb7v1
2UGSdDYEFH/Qr+j5sl5DAbALRIXTesZaV7kWgQvLS3eKIqqp769Xbxxqfl0F9kdOZzkq8j+/rGID
s/5u831MU0ih39PU7spoI1qocysdYkyCoJlN/LKj2/tcwQ8ETMAqWTZC5YzrqtTIM635a+6h24cb
8jfjHmTSKALUbTxUFyv6QOzWFBEX86T4veGpN6xO8X9R65lP9hK+zekrDrqWt0+L8axsiNyMmZ2r
2HeaY7FXCuq7PCJrLtf5AG9d6GGLs5HPRDXmwh5HYj3BSLCAsUqlbFzgNBgT1i1H06/z5/EyHnTm
sGEBq0XMSK4yrSGYln3yI2RoDHD1YkYDaSHKIubUK8JqH9Jj0TEYn9bBtoQ4OcdSgVPZtL9lrbgY
HXdDyJlkA7Qa0r7cvxxV02YWzV1iB300JX5VtNsO75Gv7hdJ6iPnKLxuTg4bDxixX+AMsS9B1PSF
j/+5OayHzLsQlsuUierDn7p7GdIaJCwcyO6L9PCL+icGpZ7Jpm2hql4K+VvEAvBQJu488ODSrWyX
f3FYuTcYRat4jjLBeSFzDzysulotMTx3IF5T5lIcLjIu6/Zvyy5SgWdZCmqU77K+75ERSPMrJ/9P
xzxzKox0n/psKR5ixjC0ihPBqymIMAlvycZvZcl32zAbwLefIuFFoMDYYmzBfLkKJQ3uCi82uiED
0MVP1j+m/sjvD3SpEevTG3S8EABhWDItwTxJVwcdp2pJP9fMVmd5q8BHrsE0H1bnOVsctbLWbKoj
kgCl4zJWBctNmurjJoI37Cqq1swilG36S++cECegv1YaJ4LlLl/Ij5cy7QX3ZmGBOm3VUmkSbnnp
qvH4rkeOEEz4UsCcwIMdphPvbd/2YcdsNHIzxEScAfDgc1Fp4DkRKgeziS1iE1MvZhVHNepSMNIn
4C8omu/onD2NZ/kdcrM7HqwM5jDq68M9gNPWPUA4EFJQnYZk7KsKL8DOkV48nomf/rIdtToKtqbd
WE9ouKc78cr8l6JdPBXCji38boue01RiLZ0txxX71VXZFlgWtKBdZpP6DUJdlppYksiuHwPAvNLq
juWCnKN48IDZd/9anfM4wgRh9KGKKdEUFe2zCW1ZdqDnL/DrZu37GIMBSClCJ/c0hWsCdkXKp/tJ
HmwIelm5DoRB7pK5MJrtRz1FpShWiXuFX1NeRM6jLIc/EdgF97nh+XmENyy78I4B037xE8OaNFUE
dKECAv6xI0Di+TB27oHex/3TdDcH5Ur7AHDse5q0BdHS+nwM673d0Ciah2CFy74m4YuhoiJrpZ2e
vgIq3pGW4FD0yQtVHw4TZeUfs42bcaX9XA2JIi4SjisJpdb4RjRXUXNsto7nukpyLyJRu2xZpUgd
wjWWfyiKoA9qguyyDgQ9n5bG7WfBp6xdkuXGlJKHffhDN8wARHESMAbpgvLhLkFhZFhveqwyc/AF
BB1/sPhAXa2hDh42X7MJUo7PFlvCE572bP8xX/pKPvFd8R2dXfaG0k2zjxXwj9HM5HkUhpS5AzE6
AQUAEEOtjNLq5qmqFBsttiZ1UzA+heT4qifj8dl+GTSSJFbMdUnPUPRrkEixOEc3R1b7T7oQx4L6
YoRWmWK8o9SX5SK909Dkkzm+hRMJcul1QPaGm6WR7qoUjX94TJ/Yf6RqDOGPJRGBtHAr+knogV/U
2wXZQnKHr2fpkd8nio7hEntV3jK80i8+d+/l5RLlzDaaxZY+MNXz7xiRIFa7zcsG531afK4PzLwP
8eBrIg+PXfJ/QfOduCfJQZb2Amr8vmx/cDcG1pt4aIt5TnESdJNXMPc0OYnZJvCALipM2t32D3MP
DcMsAdlBKQSVoiYCgpes9VjzvHt0zU1b9CSlSMArBLf/d85eZUirdg1RjBzuhxfeGEA/+Po3cKH8
5dRdEMrDq7aV6ICb2z9cL5dfEKb8jmdbv+KxwJRAgUcNPNK3ddgrShMcebjtlp93Jm7PbvF9Ei42
b8Dhqk802TXfqCYvqgT1mxv+6x25VGkYn4e9tHCRh76NpIRLebH/tA0gwx7o/hjAW80TqCaifsYl
jh3Ck4jJjyT/vLd0CbGzhJuadSkyjeStmUZEOr+TQdiZHiuD7ejC/DssNsFnqsxYvKk2dDs8a7Nv
QJ469nNGNveiUUoPIusDTSDPHcfDzC8zVmWt+97GryZVW9i7jLV/ivUND7qAAEegF5CTPkVnkDnA
8hjsSb0NJB9A4NYRgNsl5Xe0hmqPU6qnakySOyMKGQpE8IdWgOnLKsps3EPBcLmjoRDHS3YxZm8M
uX5a9LDkQAZlQ2IPWd2gWrwF+ZPLHp62faYi1rGp6i2SLSP4hsJMjOiLKe6VXBgGfzqEihE7jPMU
djrCwgYAMDzA5sdB6zzGRJYBykzuNCMuejCeYC14qX9skkE1+RnKJb4tfVqf2uFjVdRrSWYWraKN
uulbluP8iu3fzd26xk8KCV9qyyHhYJP+LdZvSh4oconr2YcWGsbC3HWsrRpqEV/jSp3LLbxez9m5
o6EhDtVEWjhb93VK9nVkgahmk6vN++CtuGwTEytK4K75Ip3tBxxOtDODuI/djvrQNL5aa+S4T4v1
OTv7nS88Fs16jZN24rLtvgGwreutSt64v+aytY9kTGxKGilYCuV8HslbH7RWBfitfRW0B7ZDJU5g
6YS0/igs+rvx8pdoka1rRtrebtEXm1FmFlvfs5y/yZTHwjaNArVMCGCBhzclxJtd6N8XhoEJxXZr
LD2U6jvkU9yXbZkPXRadPnq1Sfmi8A2ZtePepo5Syx6E/BfYhxRerlYYOoEIq51K1D2MzTEVypIT
hzHeVDH6pPJxiMPvC9nb8FyzWMxzPZMoqlHSHhxirDKUHuywZJkyvuJfxhaofKOx5VC0xD8IK3pN
ex/8yHTeqqDsWdrIvIB6LQDSRs+jae+olMCxtDImuHuEsH8O0/sNDUJZbA+NhjyTb7StUDXFa3aV
ml/rBHuLO23mKICO7F3gPPADgdvuz5UPM+6Rn3AMPWxZB9LcKIC6HWq+Sh0wGyJye5zd1CllGucm
rJI+jWZgeZucEy1WOptUJhX8yxmCdx1qkqBtQoY2q7gonjAkU3BePZNRGXGV9dH7GGUvxB9VV2j5
tOy1Ln1hqVhFGE3UDbIEFw+Z7ToJ1v16rHsw6r2bOgO7D214OSVw0mi4bKSQA29gE+zGiiBJuH1J
ldNCXhi4Y5kVk2nt8CA4yNXP6hl0k571QZzPb5eo2COEyiMwSUZEdzECQL3O6lsGKGyPlaEjyCVo
65xGZesWU45xgi2jWkKpof7JoDpiYLafG0NUzg/QZmIRxN4vWNyQVNRuMYiG4rwsoX9sXrk+Aom2
AQCZXPwwgaIsDf+kFR/IVRHbwQziQNlAuw98KSWM9TZpbdt86OgpleTJP/4YF9G0I+O4DSsojtuQ
NZtCaIemBA68KDdim8UXJ7QtIXkrkvsPkAnY19MbFCB+i/N/qWWZbxGkQGbAT3W2S0nlrYxkPe1P
miZ6L8r6yG6zJKEhyVhLxM9JByWVaTntDCeYuSe3sNHJwrRbE3CspVo8njQHDVDa5/tGQP6FB8ne
Ao4pxHAv9J4bEQwm1aTzOfuv6aAk5NLK2x5V6yOwIjDnIrqZxkwuC5mUGnOLm78Wlp7iWYUG2Gb4
RgOCwqr6ba/3/WTn0QsJ7OgQysv7PcHzjNJoSVY9LMZiKY0jEMhEO1dqXOkjsGYcHuXnCU3PvPC0
LlukWaO99Ti24E8a0bPVUrz3BAWoI4+ixLsdUdVg4ZGAXjOUBcMszj7HFUG9dQisjLRfH2EKYuzv
e2uk01ndismYNXqGhT70TQI+zeAhcBZ2B/IXbfrjZtEAZ40hLaWZ6l/9OahK1jwcBqI4XqL8ZiJ2
zY/HaRQzKbkqRri8ptsuH0klAuGJzI8hr1Ww5NSVjSJuJiOV+88XEMaYgUw3L3VAAQqoMKIq7BM3
eiSf6AzwViHcWuSOb2+zR6eYxeN62vPizO5sUSZPjnnfQ8NR25+1mlfrJ1k1jzXt9lO7qioR/URh
2yes8KDgb0hnIeVM6T9ot+DovKL2Ku0v7ps226lTdjbppso+lA5w25fIPM/6AdbrZJAxLctrrs3q
KOlujqXtvBusXrLKX70LpbUiRqRVJ0LuoR97SR70nKLfS10eYkfFBne0PI1R2FhYJFG9z9dbvEuK
vWSq85iOVi3fE0OEHo/p0XXIqMWLqC58P5BqnUJGmU3+pVXYJZkI6sT4lRlFV+uuM+WThbACw62J
eShNsTDOID3PFx91vVBAVZcKO7rrykF3uLcxIm0wRum9jU3VRW1l8J92cLoBDDZXW3Sxv8CNS8nH
uAbHH9nHcLldAhMHJh3w+cAb5tffasdwfteKvFe3iKXRbNjPHEyHgg6SPu7KCSM1iUfx9oFvmctW
b5dPtE871gEeeCZQdJhueBLVwH0f9oS4Bz+kmDjY2I6XlXYqoO5LnXKuC4D7jwA/9gLOMTeSiH5K
O/p5QQLrxd0VPaLJ6Wi0C1lFTDl1+JlHDjT/lFqn7nnjeCRKRaZvW6xKEMIBXqDtv4/78mZUTJfx
WE8BAkQqmvv6YeYdnXC6MX6LJQpXpJIUqNirlUX8YYG/t9z0g/abfOthxpkagAGWkdR7OLXw4Nzo
c0OnbiC3WupuRz5DYqK9NLiuuxNdYVk4r0iJg6QNkx1wNhcQ4qaOePL/AM0ml1jXfYZd211KvGMn
ZC5HgFSwzgS0SLknjizHB8S5odqofviRihEB5o4ZyteqYKC7JHYkOPsuWbeLTs2wBt10Ydoz+Cj0
DRACLAFDnk0yC9NE10c2FFOcrb9Y75A9nSAvEMFkCv3sVz2pBXFb7m7Xz7pefNHP6omPcqVm81+e
oE+8JKW939ArSu6dhk3U3qMdC9p3CbirLXsvzeeRGQ7APyajTdnZMXyIcnlEiCHmnFJWg/0y+WuQ
p8j5Vo20/mXw58qSKCaok1ucv7uEPyBK3GJNBIBiahPoSM265+pUdnqnfZOwd3vUKYF959sCQMkb
TGkByMzaywPZ+rxixdBg10yDurN4ZH/VUTHKfyrslqRnoKg5JMIJnRrb88XTtOFM1GiqN00npyno
zvtA4/hpozfd+zQkMnY/MHrfC0X1q6B+6+oBNia0z8ZQbq8BsX3NbeOu89eb/aLTxijMzUdCq+4X
CJ8bcL/t7chrINc5u1Gv93PjkwYFYjKyd5w8jxUsXIHrtE6bvW/Trd0nYgc8KDHny5VcNfhz23d9
pfcdp1g23bUWUkAyfQvgd8vagNKP/kYxb4I4q44AlkVUI42+yosN8gBtU1jEjWYTr02gKVdIzkY2
a5a3JB5tpTPVF8VFR17+fgpV79IuqwQZ2EMwbFtN2Mf2Fmxv+Dj9fg5yoKA1Cidtl02KqLwXb9Et
YPFzRIKac6li4Kzs1n4SsQDutWHouSu40tBHq/7PsMdUFzJjcArf1fbR8FMaXLeCLsFdmXz1VHwz
yaOjbxIApMHMUD26uIaUlxNBzUG5GAE77iJc+lcvwUy2TuLTOQk61IP0IoJ/ebbQN7z/K6Pi+SG7
zH0Uccn3t1hk6/RUSCWqqE+omU5G57eKiHozGd2c/zA9Nf6a86DccYHID+JtmVKlz6szkXMyobRe
XjAtckUZu35E56w5gXwEodDR55vsJgb/LS1eM5Gm1hVL8ChvEZg/3HijsMNxItpK9Wsuad51nMkB
kuqJGfKd3h0f1EjWYEa6qqeX5nqJp1LkBXedrQGzWm4yHN24HC5puxWsAX/bGq5RDn/XFMh4e4HB
5KFY/bBnl3WZjXSXRpHPI6ZU7nU/CYcpiIgyImkT62ESftNilkEtqGh1RXmMPDMLxT/rFOWimA+U
qYL/7VN6TyTyJZdml5oHeolcDXnjYJRydOzSeDd2uPwaST55twyWVGSsceE5GNFE0eserY3ZLNtj
SGNF4G1V23aoNsUDmWK8DmTigHACRw44cN3acEGd0gbCPR63WyAIb1pxCpX2zVa7jdk+uAqGAJP0
4PmuLA9oKCrsuQ1Tow+w7ga6tYG2MxxtaQvNN7Af2HaFjKv9bHmEMXNX0nY2HY6IGCZrZl5IrA+4
QoQalWmKsr711ylfmOlAuUEFgg0NBa34aF7c/tbxYtmoIqDSsP3JdbDd+etYZi33Qp10ARwuTk+w
Un6sGtf7NNh1jVgi9oR0G34mVTj0sbfwqDnUi8PmGei+5UrJ1jysgC5GeOggJe/KuiJmryTQgx40
yWgqKt9kfmGOcX4oLwv84OmUHV+LSpuqozBHh8pxi9yt+MEqTvTu59Irw85kwvTWWNyST8vKISve
h6UboZbuAxcmAw1utfPcYT3MbKU1QvP/MG1cjLqEFC2Fz7zTlZdpx84WV5Cpc/ikQDPE3u6m0kiA
RPkfsUTBel2O1lpa0OyWIt5IHZnr2HZX7uNL43+z0oVqRNEPMylNLl+7DArvnmFckVXAdn9d4dqP
dizog3paLlZfk6lTr70c8uDzrkxTpbNH3LoEiLf/+Gjq3b9XriIIojRxOYZGPQh/modh92BChDmg
kUtSROUAwCj1CDySAZB52fdw20Ow+eBA8guYhNbQlz3nJdEk31K61eFSKJRfPJn6G/0serZR8mdv
A9P5G77EzmsQn8q9Qiep7mLp0a5sMd6k6mlI9N2bfW+LD5uAyEfplUzTDggcBGZXrE9V/6/2swpk
FTH2ogCAOe3XznZ9pkh1cW+02NGQ2tYzNMAn9myIrz6UnGpflByxIt+qmNbDDicpBav4uiTGFaCd
DvZzUYDMTh/vDhN928U0SjZlyWzIBvLyUqxnzxf8Re2AtNZ3ZOUrf1mbzhBkUe6H9jagqEZvPc98
eLVxEbD/0lyBurVYWUvdOQouHV2Q0Cz8XSJnZeHdBAaq3B2nBVeDUBc0vAeqUHks5EbmkNRtAw/w
W9P3jQ0tUTS5EB5v7mbIFRhETeUtIDK+0XTOhRcOxynuVcTKcqVmW++lHaMuGr9WaWCstZDN3HDk
KqqH7HIYBkUrE0RMmMWJKJC1q9zD/dj0UIuPMAAdqKy3n8qe7bxdfDoohXUUDtocalpkd1sPGipk
pNrhMvKZYEfIHxgxz56uT51ZXVLcAYW+/V4Ohp9XaZ0wCurShYZvICTpKwNzP/W5gyyHpfi2zmba
JSf/a3/Jdnzm7MiW8zU+msyxpEoPetJM6EU41KHWWtDcYAafkKS4i9QgTkzArPRlViHswHsiT2qb
Frumy24N4BTL7BNXfLQEQ/LXxCeT6Wi+05b1oa0QBbe8CuA6PGxLfbra/MFbf8Euw+wtq6PNMnrG
B4YwE4e4bj/QdsGG4sA+gf5kglaLOSSpYXtTi7f0S+Q3suNKcmJUCoqGtszDa2117yRye+NCwNQI
eIFFrRf1xa/220/yL++8pGIXuthnWYyhJsJmhj0qvjWExFdsITsqyovUYTzcpX3DXtL8bANzoLd2
RiEew9x4mwvZNwbBKwaUXZyrv/V+gRcQaJPcTuoUXqP5aJ9YMdIKMnxav9xyH+NZXA5WmD8ajxzd
34+bxc8VTnJ+gncwXXJaQSLvKrpZCbSLCCexEK1lZcD8xUodOOGaP9C2TAfIJa/8HbtyTvNzZuQg
xcVqMvcua1vVvDr39QVCLeCByPGkbPsBLGRyJdBelnC/QSCzxfGpUOgINHZ6/bTPj/dIj7iyDByb
ycMmY9bkf1Bu2IFibljlGt4vYLsMUdNyJQr9KlT8vWKQT3Z4hss/u3StCFqe/7p46eGJJtoxwcwO
52q6Y4RqEG7kgLH3GT3tRDRiaJ8Y7uOkxb0Mo0f6BiafeIRKRdbaSWRazMrbLskNKjWIpObDpFWs
mqrJRtboA8AJLNR3FIGD3co73DrflZfLUqo0k+ddsHhG0V5KdaS/SsT5cvVaYaZ3EBV+u9wdRtrD
vPw8QnGGpqmBbRTGQU68qr7mEmK93ZorUIpfUAG121XqUVpcGmbe0Km9NDo2XlXQAqmE8e4RE9bY
+HiT3rA6jn5KMONc/PKKXiq1uysMeEFqPxtWKodAd36M5g5XsPLbvyd4TecVUhqPTezOjIDTyByq
2rp73xmxhaQsUsUmiOjHd9bVTq4bp9h575J8LWN/Jylos06y6NEcArevCdvBiIT4rBqsuQUgoZEl
AJxD0KQmIOE2ng1IMMCXZmboA1rlTFdID5siKO8DtVARjIzRKu5mjrGLh3lXWfg3xYp9q6Frk26q
7/IRKj8wBA4aGCvumGLzLKtMm9zq+IK/HM+WiShkxe+R+dgeYI32mYsMGp7CNEwlqCM+BFzzoFHy
lF4OL5yLHpx/zrZeSFaEbc8ewEH6FXti5kpHb4y5UTJ8LDtRWjzDbp2q1+YVzXkpIosPSVXprmLV
j5WZ2gELIqUpE0tisHUleq41zdg6f/Qx+moZ9IRpEIYFZCDQ3I/L/+CA/FFK9+kEiv/IK51rZ8oF
ZnZpbUbO0z6gW+6/0AnYxBTyHcGwzUYpW86dNWefcifTf+w4maL3SXhc5c9tqmdKxrc0VcbYTzIz
z2UupcmNNp6/tv/06zUd5CXCh63ilv4CRRThjM9QOeYS0NLUkeSZ/lUkoW+17N+9fk7hph3qAXUC
2BC1IvZhIWUq1l1fx4vS+vynwEWDB/GK8O8Ho0vymCcna05xbdvFoWh4BMeAwTNKO1c5z8a1X4vH
MLP/29tdb0U7KgTSrZ5UDFKiy+QSAGj+WfbSNtuUkNSgkV2iaLWlKVi97JaQThWsEvFfWjc9CI/5
RKLitokJJai8n/5lAnl7W+eqjgkjaaBxMBbj8coEaeNrP1XU9K2UXQYUi/keBbe+7d177v7NYJBZ
2Ri95CbXyyw7GNV6O4S+Fal6un/HH8ASuTP4DFeLB2I8Cn5miVDGwE/2LIqkLolnrgjlTZ713xI5
Z8HqwCWyhdQnGevI7Rt8nlw+GOIKzGZt6F/w1MaBvcckIX5KmofICKScrx6dkvQsxJpTxo0xgBjY
kocozUYtasMDUwemvvHOQh84Hcn5fF7JLUSVCjSBex+q6bn4DwNg2M7sy23yiDXz/Zb3TOf3zDEH
+93tgprXM4CpaKd6fLsH9dwKsLSRLmdYxExh2bATXlvv/mJfl6jTF2MSv/npn3HQzPQAzHBTC/BX
KdFUTyNqFdeV9Vv839/LimntjLfcerZJRPI9orIxirQlnzHMuvTYr6pb7WMRtDxZt+iTOcgoIIHZ
sXnrfXmNmOo+VqpQD7YJskUhOhUkCDEIgEwsXNCooua3SbwnoxOd2OoWCfrfblnvEmESl/XMfPCH
SvhakaVcSjk5kHPsrFDwQSrhuwS5g0ldQzSVq81VgqALjrKuB5/HmhGxl+4271xzmHSeQ8/Nmo+F
LEFu0iolykyQpPEVxYgdGkbBrx4057BdRvERxgfr9m9cR+hSMjgmMRp0YI12dN+GpadfP7Z96KAH
o6U/xCDwVzxyEgfgCrGSKAzDtkodSWVFDvv0AHA3SNuEUn+hWBSfIHtTxp6V/hRZSsrcmg0avrsf
AVDGSfWooseR34prhf0STHOwfBKH42MUicYkS5ATQh0OTNo8FQqd1jfv43ref6QGZE7KnwxCbHN/
vHKqV+aRwcNPiWusf0ipe88IvJq2eS4vhKsPO7Dheg/BuZzHmlxmica+5GVLyCL9MPXCYPrmkHIB
UqYddLZN43nIO6bKCUTSxxkDDJstuurdPnqvfkp8bRGkyBULotBagMa4jDdxJLgxcRYWWlEe6ULZ
/95Qr8AmJzni7ThSo9ukQvCoqpKQPpYN+GuUHQjSkp6p48hg4kJd0dVCOR+cCYHbbScx4hugASJd
XggcsaSw1UZFrXbUHxfbWl94lI0VMDPBZcxNj7zC86bvRq/0DlveGWaH4HEqc8/3R69fYI8YRiQh
4dhN/NXRihi1RaLKLTci5liUkr4C4QE8UhJGiK3FGSj17Yfh1AH23jsBTtZDguBj2pgpKeiyMVNS
ohRqVU7Vcgeyfxf1Augbf++HRsl8eryyCA3TaATscJMQc2+bzgDXDIcM8D3qoqXVRsOdYw4QhCAi
e4S59NSnNr55dyu4zwbbfinadj7oCTDm+DPtAHzp931rrDewOh68f1/hPpRfR9OJj2YcWDr+1lmB
Detm/6iODjag7E7YF15kDH6Ga4Re6/6fab4J4FnUyXR4Vc8jK1pKtP8DbSjPQwAOVIwSO1DF7zCp
kfanFab0XXTMaBrS4d5tdBYnA2mGiy9786ZHNRfeQfHdnSZZ+UO3wSx1ctTBWuaq5KtTVivnG1lR
qRJOjgIX2SwQw6Rj7xGNsyqEN4TQ1Hqngj3pIyOsFW50kNxuxbcqu42MO5Akk9cpLQi3iFtGcw9j
9/8viJlm3gMgmyC8wbDf0P2Lh10TBE7r/90Yar5Y10Or+zj4WppoxO0GtQZq1GaTBuGCuPZGSH2+
ANePYfNuJAtOMbzpT+x3tCjCDhfgg6QqVpG+0mA7mzrYWrgRSyqZ1nrUzdnSQ/mjNbt1AgtpgTVP
5eJKztcyXL7OyW9d3mIxxe+7YYENHnQx7fqa3seuPmuVi2JDxDp4dAXc7AvEDJBe60OOKpAGYEFi
ZQmLSqsBMNNjWQUC7j/XbzCTtDYKQDej8jfwU5XVSVD/ce2N8/YgNSPlAOU1f7S0HFYo0HY6Ruxw
7HSg69QOXtMEkmWBHPZp84Mjp0pUsqlJceA/42a5xJE/stlstqdL/yjBZqaq2mLDURIQ9eDQy9jJ
v170XMTe7DsnT+1yMEIswoIW8czSRuIw9ADUvJzTpWzt8HGIKlR11+F3ygKwDdIuEBvedl4lvo7R
v//ocXInUNqIQAO2Ns/NQcPWKiP9vCao7GE/XA2EC+dmQeI5OTw4OmCn4HcbainFVlT9SH4X27mL
j3DB6POu7G8A5zOS8JM6DyzB1FzXOLWdlg1Zyxjiig4rzfLRjUd7FWhTjEsQCas7APr/VBbBs6By
e6Sq6jGHzOsCAJH2/8HyEQKg0mHZ0ErgmIYz4L3gHg/WOUidWOd5uarp5F2e6H576YJuOpzFJHoO
2eKnTIfHOQH/bVtLaG2v/Ex94yJ9/a6smDSmBrmPc6hXRj2nHS/jzfljjVsnDq1gpLnEYmv/rrAc
STwi7n8rcUDrNKzfI3dW+yteOSajcomsEjhoeZhPDsoBdL72e1V+6TjP3t9TXwlXuCuMGH/cll6g
+/KHVST4z0/ecHitpj/p0EgJ3nPRtRLm4sHHGewl+r6+Udotx5jrHkAhSWqS5VEP2C2W8og/lsFM
/2kn/e6eaahp+VSeW4RjvmaFa1cYYEcWPLWm3MbTsZa+Lk2Dd4TAYJh/hSJXbkhOSJD/aCRiZ6el
bnPoaGIObAG5KkhD8EipDw3kXUub8AKXXvDmQNQD2tuESDeXx2AODUuJMYvEY+lA/LEoW8NLuaX+
8T3OAOL9SzQZjk4N0BvT/cRN139pcfiOBqFxqSuZYkAMquCqyntHKLP7yWyckQZHDnQNIYwUGAdC
48SpYwZghcfRueILbWNoMhbXZhro/woAU8qZ0+DWYTP68Y1LdAXCVa2sDAj/k8ejIjCN9TT50oTz
GhtsLlICrLpcGGeQ6lod8Vv7+l5dX4nJLDMwg86Sb0Pc9tQPDP9k5zwCW3uyR14IROKgF90ZnhMp
3yJnfIc3RD9UHECufU8MrPIOuWQGGWMokrUPuyiWdxgzPK2gDPGUs6CP/qJvpCOXdpMpvknLFy/q
C++s73Jz1QvyMnX5KPgxxqUybMYnT6CnHlYRONyLn6fLETyRiEW+PVEAnlxd5viyeB76ZHYV397i
D3JLjweLaPd2JpBHav1JTH9UrKVfdbVTJn6KSOFq3ZT8eqLpginOuRZfidkeD022yjpl8iA7r1PU
zRTu4kowGUjllOXOdhinEAILjTVw/hBz7VZ1CS+n5xe0D6MzCcAASOA0tLx/acJKOfqSIpJIWV4t
pwFBaNqxWM3IVzBJ39qKVw4t2Sp5Xpv+FC8v/O2PeJ0XoHaIlKniBsl10CQWoMNMLHWopdqqBA42
0hLUbMT3lkiEFz0JZRwwjZND9Nl5ZWMAoItGcy/Fj2KFke0PWsFE2wxxpIqRf5daL6fmihuJRvGk
iiwlk2j4BTIRvQ5MWzWI9bVh5HTSgW9jupJtlswOjoccGzNW0q0E7SG6BXpqwxgzC0EcpMfozUsq
f8EK1JycdoFYSsTB8rB7RiLayhi1lXPbm5xd+F7DWV16bFbHDBVk0kRLjWaeO/EMI04VvjZElX63
Q+5rqHqSfrT4iNfcCDpm6KNSRDWa9anWaJWB8R5sLUCBfWUS5p9HJoyI4TyoY8CFJo6PEBCnVGPu
K+QeQo8eGd3XSyrO+FwGwPDivrAV1iuaZt8rCZJoCM9N9ao8WYcIh2u0iXHKqbGL6fUoPoyLfRaz
vnht8QARijjHvgTvnSUPAzYqL7TUy0FGmoHkKkPyNhJEXO5e1jCS3y/NEvHsMU9x9t+p/zZIM1v3
pzB7djVaOXfQTWBL2zSLsl/LSPH4S7L3jJXeHCKSTVzCFVF32aE0Jt3l/VklSQGf0E3cGw1OzWFP
zix0XkGiojFPsg5+lS6T+nyPgA9RMSISykYAH0mPfWYwqd9Pp3Y9655xLa+uVefQd8dnkG1kcZoi
9zmvr5xvOWaW07CV0nGMcwEShEKvtUdxBXiijVkG2wzr2e1E1wnrxSfnDDA24QQY56gbnPvAmqqd
HKGlcVwc2t2afLA3fS8A2V/BEmyH3U2L57gaDvsJo2HBXwjf0wu3LDEc68AFJs92hHpc8hIWQpLe
sNUGC0j3q6CA8V5PdBOoA0ybRMcnR2Nc6+dbgKiQKgGAl+mivlWZ7DCZYgyfVAsg7O1XxiK7WVmn
fmYwBTtjmtNJE5Itub+v9EfRcebwsuzPYT8iC/UrG7Nnfb5vOfL6+sSDU68GgOptORO8NULsFnwN
07lyzxMyYiOrYCuImdFq8fUHLLOx6+4BsVKIxWFDB1czDywNei03Baz1mHjGhh1af0hheFbWMWoV
JZzzOxV34ybUs/5tfAk1AmnELE7X2bz5H4JvE8THK2T4pLrSpSq1ZQHhH6r6yn9GPpQRw2BRuQIM
iFQ9eI/d4q5pSkjQ42eGpT13rPhxHoePuF4cvxXTwTmTJJthIRxbLFgyuA68AxXQIDxbxphH6HSS
mllVnN5PjIyTErPnUBQoKzYCfZiFGLaFYx5R0vpvIorqF0z+W1ZSJw9Xs+zPQ7WoBDO+1TYInDCT
aheBW7FciWX7bjNyy4Kh9b3HMv9aWljkRhoH63aMaetWEJ+oPxoe0/ilUbR85WuGchMJNMg6WLH/
SPDvcEiwPsyNXzwQEd4MHSAPw5BfHbGD3x+uPDeVPj/FLgHQRnLYpqVX/CBl2AMhZYuijQwkyU0p
f1TBe8FMkENpT3ik2Dx74z+aZBUNGEZSZK8Yq5Wsn+yjLtg6JvUYUaBhFo+5Ecv3AGwB/R2ykZ00
Q8JQRlJbFyuIkHfHDuY4aVCO56kE0WMNsQqpBlO9xVOxVx9xg9iaIiJmKQV7dOEmvOXrH2xuSQ3x
OBXeGVwbSsHdDAvOUSv6aNKV+X6nxGxAJ0unIqGLJZ+KyWdcY77ZOOxlBTV6B1FXyXki+781XsqY
X8w0v7BDzR5Vy9xxne95m/6hGlmXCrmf0XBO0/ZbyFgHDO1/eSSI1URg3weYz9tljyqJw5SfWYaz
TYobDQn9xM5yne1yILl6acoe/7QZqBgqmW0b6VFMy7isA/tqMi8aCqYbtBMOVsBfPwpSfSf1UiVH
J3dwJDGJ9TVeUVlIKCjDynkRfdF0W281S+5ed94/JieGW2apTJCgUblEqYGN5Bv20F3jjKBSKrGl
BWvGpb9oAUTv4OBdzGj6Y+tLk/xdTeUhTcnMdK7NA83TgJ7rYdPRdrvEvPPkb4lH9c3+GC2EFzQ2
pdALdF/q0hiHt/zeNV1WrV6O5pwZvGKocKOnmCInoGu4p3JSvJj401b41aNnLwn1pAIT2n4QN1kM
BY1i4ynIa7YSTtTH5m/A8UBPiAjLAXjqQAGYYafpScllYdnIvTICz8UXw/zYL5rG3ErwFH1ZnGjc
hokYAbbHyTKqSSnVMywmoF+dWl/aVBP6SBKMn824BN1eWNoXA478+qa+boj/YysbHdsckrSR6tg8
ODHZaHju3bvG356Wnw36CkVS+CnomG7lGCuTvMiOBqd+iAxdQW4IwUKnVkj8Rj/7O14QNYXdEBA8
u76CNd9Gwv0er8RqJB3b4GxUUAZF5njORMvobRzF1FDX/1Ri53uh5D3NaJu7YpDME15RxPLBHYtm
3mctB71lh/DrwAsFrebMI0q3ua2pPiUsgxIcln0j3o4k7gdBs12226q679qhSgU5+ZLz0YjNZ/ZG
+tHzBD0PPBD+K7GLF1Q1FLG5TljbvG9LBo53wSUd0D2aV9RZTJVoE/HcBbBRGOsxim7KPrqGrIY7
DRU56iZ/wvuehnX7yzqOzTy5xyOJudvry2BtnxUgqN4+V6zhb7hXjE9PaxBoObSkuqwfYjXQlfHr
1b4riDJ7V4lhLqhn1EV9dtLAd6doqQyql/2HFM+iB21hFFt7E6GTlrR2KjygVa/QggGzcR7QMkPo
u1zuerhYxfkcLxA5ujGoyiXEYZ8wLU4pAsYbZs0uMGuBgnIG4pVBZ2KeGGj6l0UCiIwax1RLjl3Y
SpZKX4+/vP7VwO4Mw0OAm/DFpd/XFcYZIt6UHDLzIeOyW1vFp38XDpSaphcXrp2GD/WxSJ9QRqbL
dKFdyvd6CmF8ySWpfBWgdI1SBQHI+F9xFSYnZj3qjfvjSzJlB4I/1Om3a+zMWhgMQyMijQA+sU9R
pX7HH4MATqqP06yUUgx6SO9221cCsYRzuoXjQOr9ljY5AmcoQ9O5P5DBnhAh96GYpymkBhxXfo+z
tSRcrK6wVBgnCl09H0I5bnRYKpCIKjk49SgpNa4s1+Zgtzf/6nU5NQIjGXu+asDA8FyPzLn+Bvyc
UfJ+2zJXIJQC05RIQeFwDpv6rK93+Bo1ArxZIakmKSlluvFN/gW5lNRZsLNvfl/uTX5wgGeyzFJd
5Bwl/BjyKikp2RMFgnDYq2Fdd2GOhXi7PCaN4bHAkZZCAnbhkpgvMbnXxxDGoZQa3IciE1sZRGYJ
7mBkKr4Xz287Hi4XEd2rzgZ+wB9mjQcwuhcrm9gpgDAis0AX9l6jNah9H1UDXMR+7+5Dp1cexakW
r4GYoZOE3EYSUM8FvBfQv6KDdnytZaNj8DxBIeVeYTJs+F+koXrb/OeWTG3kDtqBZDoNVRzvpuI4
OKGM81PWH8evVSIrmWIeVN8ilyanwUL6enptD4Olix4rFgda5n47TKfTlxMqrGev5Qx1aYjv6x7t
20kGo4cvGD1SIEBRXPQjcIqk6mUGk/g9zqJRXirEPUcR2t2syrL9dSYCooMz1Jway2EL2fdr2bDJ
bxMDnjv/fQr62HTlStM8EIdR8IBPzDIzUrT0+K4BfaPj78942LU4GdEGXVOMDAQuAYTXPjZ+gZC7
LPNFkwTNQuE4ePFtMcG+iuHtZBH+IFFHz7TEDvRAlu5RRnyJisXiMcy3QmwKhXDxDFEOwctmwl7l
qIbElvx8ULiiJOZ8BEAhj1wZ+5QT3Ht0w+swt4cf6mEMfmhlkRBGovQMlauiCxej0wh3hobflp//
L5+ALCinTi5HYV6iuLqI1iN/GKzKXyVVJDYVJdC5THKs0xvPShcSdeJDMgWj4wj320VsNLr/aIgD
VPRr1c5YotJuSrnR6rLiBURDuV45TziZHzeFUnD7JLR+zJjwvu0eCjRg+jH2hijbwzIqpKjXrpiH
RcK7ZB+t0DUMl4GwNEFRk+cMJkZyKX5ceuh7HL/5zh+dQ6r7cvZDvNYiBXziePhb0h8++1NoDZ4m
cj81/OUt2etx1A5XrK1kgEgY8S8podvfQ3ovEb2iFvNJkB3cK/+TyioXnn6L9Gao2MzzxgXiSCNc
WCYRilgurXCNAY05xW7KaajjCNOLgJpnskcoPCCzG3gPIkaBmyepwVv94dEmY+RCnX5wsoLM/n4E
LXYvGy+2EMdbS2LIa09ojMwLFq9RVkFu1XMGOoyoUzCefE1WUhdeyzHCVod6UH4U6hdT3ZKnw3yQ
gDHLiDJKL1oZ72wouZB4j4+F0jsekCyzN9Xov/te4jGNzg8xduSbS2Qxo4d48/8+esKlvwqyruBC
ytaD6pgaXm17JSCsgHu+rFaMBSJcqJXyj45AC0GQ7wzE6SnTtc2EwPzbj1/1j4OyepanpsCxrcqZ
LusUPMWESuaLpZVK44C/PPt/AFurGftQceVbUzqo5Ey0erG9WYKmV2cNWIEuJv7xh8XlWLqa/Mp/
bf5DLtVfvUeREMhL4JvO08ipGGU4eEQOfJs6pC8oX2/3KCEhxIzKrS/bm9AJgdWN2NjeRelYJ6Az
T0Ei0Dzm71inlnLxTOYSYeYEdVgvPlSPxNA0ZIrDUFQbWObL9z4Gqi7p38UG0RlcAy4Q79PX9Bdr
E8O3SL6XF7fMiYrmB+lLtx4CIbHmKIg6cSrRX9nzqgJf8sQoSJMhczz77Uicbgrsr+SYLI6VHvaR
YZq6wKO6jQeawkPb1i1S2BJYdUJwKNVXERJGcnk33Elen+5v0MrZHB4LLQnXWrbmBG4Syy/Ovyx6
4vNydWctwQrcJKBmlrVRvdcz/mfqBfYx8MCzAWdjing081momB7lq6yKgkqDOo7c/dhcn1BHn+KG
YxGeV7sUewT8JuSWPPbA41C5aMq/mOp4FvsREyK3E1qKjNk+AdAToZmN0RVZrPzS+a1/YuaEnLM3
MnmMP41hLRmxS6raJaE+h+bXi1iv/3GdI+g4Ze1VwSON8iw6cs7M7wJZwL6SrhQgEQ/0hsU55dW7
3VHZSuiS59koaihgvMUyrlnxseBFQCoJC8j/7ImNENWC5Av2Sh7wc0fVJ/nq0J+sQf206Mmgrle+
5yFCnuVVSKJC1+EfgoWiqB4pnevZ6xsdTWFwQpobu5WnLS8qr2tbPHBsLLDjWP+KlTpw5tYhaEcg
zKlhOB2n1oYuEPQY8U/rVTfkPTKDvsx6EHAlvN1pxG6jQGaSZVmAhMLFLPjQkKPAUJipX0o66lTG
Amox4CGrINXASOQ+sIhvsyXyKaKyit2uF6pcNatmtQbA95muF/6tfQLPKb5fqp4+GXcdOkK7uBa0
f1E89Bs2ZtXJx2M2xBAnz9iQmn0pJvRZ1FYHSY3W79GIGL8XFUQhC0nMyJqLPjfKkMSlXsphyRAh
eEeM7Uqj9c8KGGl7I1CU7SCsw8pkDhGDGRtVGHXTIG5umKv6u8dkr0nbGprSdfuVhU2FCBjww9U2
FEQMZBUVzzig/XBnjb812GD74J1AVGV106peHyeIghxeJUudIlWWASllc00gvn8x359df0lqKoH2
qQ/UvzpzmDUB5hevqZwhl+MNtocyGKdjEcJ4/j0Kdz4bElXEEUkyPy/XrxhZQS9p0cUv1TTWkMhY
aIOmx+mu0KWiFZs0+AKM3UFbS1kjc9ZWy2x+PZ0hRyQD4jUaEoiG+lQLJqSKdOrDawQ5k2GNZta7
mpUcR+kbftc5EAHTF8sFmi42+3nDgjJ8S8QM1fuapOZ2/jgKhBIWkNYfLjcpcCKrHy35OTzS6bdh
vnPEZSjoCyCfsxkNDVNDNUAfc1jzBv0BL24NGLJ5Kor8zTimSlZD5UqzqzL7KSVN9w5NQ9+ofO0S
BDp2XsXweK7eIpS0ISmmkQ0+QTDXjCsm61dNBkUHp/coXSO3ouniuZDGcyR84inXVAQ0DTZUTqod
K/H2xypy7b42lXN0tmiDwVOTHdSKlm8QZF1H7HQF6xKIueoWt4yIoPuifBFW8NUwx8QheY4qd3ru
+9icXtQi3A5x48aVw9OhyIpR0VhZEuYNt/9pmY9CRq6bXlyEMXYMJWNulKnJ9T4Ymex7ZKjA8YTu
H6+NnBks0D0Gob28VlZjpzqVvWn9CJsm5wiy0TSbdQQhNOkF8Xguh6pf4MshmE4Bkwb44aw8azBy
Tih5lYuozDg/SM3BLIvDHLOBEd79+vRKddhAD/bZy1icq+becVMJUH93i1yzVGHDyLBB0P0NHORK
HzjR/DGT0hjEj96iJS6fptOCiHNcJty91MgeTiKK6zcsad43vqTufcb2Fqs/WTYMMpecx4fE16q3
/HHW2NukoGm/VEAoMP/wQSGauOkT1OYWUBJUcUP8AzVK81wo2Aa9r1LoMe9os1bHIhHTKsXE107p
fCaGSe8NyNZsRR2VldPuC+aeTSkSyKN0boXnAD3Q5GpdLevTkoWD4feqJRPKoLyJLbKqABpLCQU3
1QDQTpwVBdbU5LxIDeV6qesw9rf9AYv2hZNJIx0xXHrO1uts0SHpNJhkKB/X/MtzMtrD41io3ptc
wp5dFU/yXAzL6WxK3ofgqoowh3S7xeOQR2Zq1z1rN7DRMWkQ2UzGGnoj+jSJFIodrgSr1uEreeqi
dNDPtbbQYA69aTcvkXIsSsY8vMmwlusXZSzeKWjeV5tPwKgOSTUdKWrJ59P5wj4daRftkyXlLA9X
u7CFpIn8ebm5iwr2DxFO5AIiy0zqnuZkIieXdhThrnM/ZRJG1v9QDPUSELslFn1s97g0V4+6pvE9
LjGRkghiz1ghkSk/iGSXHgodqUwjzxTSX7Oel2Mn3yP8+a2WHDtnAzWfj6FF8YfKEznznRTvP2eJ
cUCyHoisc63X2ooPdZ1jV0/vgPoVYWl3Fsyu9dIqxbONwpr5+/iIvJp8dkt3UxiUNnE6gLwZWY6s
QRpxu+9Hmxx4K9VOgwg1yXV9M04uo3FKatE2e7+5emBjrG6EzaGpWOOrY9kSxUzmumHY/CMcFT07
FTATjA5PII8snAvI40uSBBxkCuViz5X3d7BcHtpXyp4qovTGQVPj2Vebf0LLmzNOHBWPLp5q55ES
TxVjUdx2D2BN/vrIIfj3Otkx6itopK5ydaK6YQz/lNfEbHLw5TGRcE27QngsTvWs2wAIKswue//e
F/ZLPxSAY7mKXubXEoDttjwFfSa669rpzCqaBaxcK+zprVRoUSG0IsXV9fSo8v+78rOid2GoDCAe
8+BWm553T7Eww3rmritxED1KgG63NcdzVczTSXW5hgp+IqpIemOun4lRNGJ4cE7xn7Z1cnzUyC7e
MtGkKKkEwMldjFngC7cOyANIss4tBmtQt0WSOfyOmsqpB6tKkzcFScmS7B19so8RzCUuyp8PjRai
CrJ3WfPqfzjhcyX0Kh+KaeywOTrG/ml9UOdLtS+vd8DQEwrfBNpt05D9Tefy7U9YHEAw+ExQl4tb
taSNuIsTJA+jQxKUsPO6OeFZuUhJfp23+suvalUHbymn4t2o6QNXM3gGNxqz09WUJj8h2snAXg8M
dm3qu4NFApbeKKBaw0cOPHPLH8wGxL7ac7JXxlXClMI/tWlIi4QVEApELaDFMtr3tue/G+Y2ZTHI
Xdb+jjyeRqZdKwJ8h81SIK+80WiCoOHIQnGCO+Nd2K4XUEQ4wDTg0hm/W7hc0ry9W3Gpu/7kd3QN
EcEPxJtaPht8l6ejMyYOtSyBTNeoiklMUPJeIddiZxmlDsA4tfPjAuVSGidw9fxj7+Ec7GopE958
zM84FMP3cLnbJTHmYH/NP/y9quTbMRY44hn6yAFpA+eGM6NIfs8GPz58epwrRvHXUtM3THGB+gQ7
YXr8AlNOqIWJJNdhS3xNzIG8H/QdjtT1w/dNBN5627q6Y6bJU6iwtrnqtghABt+s07SMP7HvrIWg
Za85vXCYtlJZu/MtvmicqjWZX8AFui6Qi2V9rvNbdRAcEsaPZlIpp3aH5pvI+XH7Fp7KP27287B5
y8N1xRiD9tqPdPFatXIMUojohKxB9L4TtqNrG1jkeaDzYf/iiYj1oEbTZLxCG7x+Tb7a+W6jd3ah
K2ajhYnBjuUPpwuyy5mcbA9VTn/cTWcYEsBU1sxuttzgZHPFsKhlsiaPSA+8ROKjNL+rxMbzaN1C
hZ7kMLzWgr8/s2izla4+hPHyxSydcpaRBPPg9ZY4QPNqB4xn4T01raGVkhlbxCkXD2yK4C1Hk8Q5
DCdavonfMDnQclRKdTeomm+nXopG0aMU1UbE23wF7dX/x7vvomUtsT7WVx1fAAMYnaZtMlXCFZnE
+uPivvMM58OX48dl8NJwcHYHYLNHxHLQjOP143BfLaBG81r7VfcqzqLCsmxtESndLq9Wgl3O+B2J
Ijjon2mcGi2HGcJyf36xWe8JLtQnjMnE1Pizs4tFQdAooC0ywuzN7WsoGTUWt72sAAkTJZcWEHFs
B1HDVlD2yZU8o5Df3usi93GulmTr1xZUAuaNmkFyfp0inrEyykefjoEooQVHrgrv45Ejpj7d0tZw
YB0wILMQ6Ii5WJ53Mq2PR1IIxByt5FRlVIm7DEnaL6MCIOWGcU0bumWJr9yetFMcpgWyyNJHNFRI
ZRTJKgZrmF2KZtrWyZG3Ez8Y23JP7OfJErUd8uNbfNwtGZqgzs+/UEiIrxLYCuydtyxMcspDZIO2
2bFjn2cghOQAM4AZgMMpfpdamOsD8NQOVW4hitAc+0dBKiOa2iwPh0ERpPmTs+O62TAFINKZXsnI
5C8lXFnpuERNvH9ez0rXfxZtJyqAvSTnzdO2hoTe1PP3Orh1LJFeAN12ZejcNPoVs0pWXcf8TvWy
R9fJf1Yf34xQHM/AensnnLnV6VJsoqv/X5iSkh30aWqX7R7QgLGF9VIHpo0Xeh7EeV6LCQLufRjE
v4CYowPr7hNs5W/4pHBXG0wGt2/MqR9YLvAg08S9KZZdVwSX55H8UaJ4gC6VOnVskhNnFHBeBH1I
mZ3T7ZPReUGZ9ng59NQDvniub5Em8Mh+zdPLsiq/QD+A4LDy8gSmMQo7rLrv6XJnwhI2PXGJC3NL
sMUmogdXXk5xuYXYhYeFHmfd01gxwZLHEO1444moPEgPkeBJEeOPx63cVjYVG9b88UGuXel0dRER
Fd6BjQ00Ls1PhRfQfV9LsKE4H4RxObdkOwLah5x9QaVGXc3ZBvG6Tv1rTf15yYeXK3Fe8L1eo6iW
Ur6AL8gg6VNy3746UDtDv8lufpjHGfyM/cny+iGM6w8gALf5YhammjnLLsyaeIIELU9kBMUhIRgw
LYrfD+S6i3zYueCFDg6WD2Y1VQ7GxOEV5Xi8UBpLJ2B1I/fnXDnitNr+XIPlMnHsVM3AG9AP0DPA
wFeukjS1D2tGBghM4Z9M8vBUFnQSkRKz2QHupDMLjEHXNIBsnCpGfkCKGzj3+xtlCPENXChg1/9h
Nk508g+PPWCyxHNL0hvYYYrJS/OR4wWlUSBsEBXar4fsRYSXfyuX1WBRHP8cQo4x1Ibck80scn1q
oUuTqyVaFfwTariGbbMO7eBSKtHhZVpjl+QfTQvZenmXPGfnNU/EHSzYBfBvZAHq8RYm7hgLOld4
V8BC2+M3rf27KsBDJ5//AG/7UduS4XAWOZatV1lKgvI15SFP4myuRa+UnSVkGMc6XU725+uo0bFY
NfJM3aaK4G5I0t8RoV8gBzYKqAL8uISXPxjVcQTdtGdZY/kmtrDXXNOZZMf+bMJ9/EPj6cCTBZR/
htSLPbyI8YrwEzGZ4ehTDaWv89HUMaKHZir7JdTyVqzVMY5qScY9zfYDwZRkTY6Ct+VjaDghKw9s
gSCdcyCCOqp31szMDbYMJSmUeWFajO31PmWQuIp4bzroAIQ8ZXf13C7GfTHwPAzrxgDcEsQdG2KN
bosxKVHOyt16/0Rz/DOx4s84Eb9Mk9YC7DpyHNhgUHviWO0A/m6jR/zvc+sj1V6fn4ifv3yyW2qq
WFPHFUyu1pwY2BdpT3IzSNsUdXSdeYwHLIqNgOoD1rb6eQyf2khhWSmk3goh/yo1eR9cXjmi0uK0
L/kah6uNzsW4p8Mi4X1lNhjf6ilvg06RNGGjZ7xBGKIssf1btm0CtCKaayNbdfl9QlzxNHTi2YeL
LgJsQX7LwAqu8SST5cAUyrY7iqnczMYR7b5ygJSdKbIpoNV8VlUy4PPIR/DwySw4CkD9+L7pDqvZ
VZkbfdZcdViWtuh47UykRhUtraM1i4gjb88PPzab0hXJ6+SoMwc6rynMYsNwKrnNfWNRnpNcy3qM
VU/4j96HAVU2VZ1YqOb3pRF+VWr08gB4msHYhdTqUkEgN8lkVLn9D+sAyHPsdc1PtiyreHyOjjqg
RrxdBe0Fex+C6emJq9Y9/QALGzu8Cr4X9vYO/SJgJ/21CRWum4T9ma0xJtnECBg3z6+C87dM14JL
uhbtjM3y76IXTUCFSY6t+mrzXfEJjMBpp3MVszQrsODjQSiVCZhYIQ43jKAjMyKM7G8eQPFCWMnH
UP6HjyEO4cWt+1fS8DtvbijAVGLxM9rbHTR19V5fNj80nOrUKZNBr4D9YCG2e9uFnPI4ACpH+FBF
AtpFtuEBLFRvA/EMeb1abadBvyPY7D2PYqXT9A4AqYA59zU56wLdtHwauDNgSXIkU7bcJGqks8Ht
wtdg56JhpBUMXndfuvKL0Ru1KpQz3MpAKmP2CSbYwRSCpNIfyLk+tuCmkMGkjMQl5faq5leUxrHU
HWJ8L8l4NQGg+ICUpKiLetyTPX2nyK7UBb6fZLS6qKEqcZNkMDaEXwqOMMyZGE0eDu6ztIrkL7i5
5/c2UOd0An3PvhVTm6J8xMFMwKsRhx5AFT+fDYm4HKHC4Azx5xOrmHww4meMb+7KxZzbo5DiNWyt
4Fl1IjfmTYJ/ozi59UKvMHOaIo6EIelb7wNee1kJWgW93IZtz3kbjsJaVJg+TSOISgbyyORNDQki
RIw5c31aNae02vZOZgPlPEJtDLOatyvk0KKa80Th9Vgll2LrPAxm7eOUDVPJOx6qGqTTglMSYxoR
04JyM+1rbm0e2a2QdVIJBQYbdgjNsLBRRwaDAG0JxVPczU0P20MlZhtfaoujNccaAHNdjiDvKGyE
2qd5DqCEVAlOo4tU1maTJ9n2oKlzJjdOJnu5xkC8trpWMKruHAtorqiYBiRiY9xU+TO/RzqGPb7u
1RWrxqfR6Lqm7RrF1UFdCbu8bjIPH/xlQnZhvoWpvmAAmvp0ho7Qn4ehILWV3o4fxY+iTqHv4HMt
DeUSPX0vBSZl/DLflLTTteYQUdZQeEszLxtivPxRO37Jk/tAdTtOjj8hxLNoSkpWP7k0Mxyy5sjE
k8/XpHgZCQ+1y7dGGoIynztncGQ8+7CAgYrynbaPKlKkB1Rsoav9ZxqLcC8In73wHYxfjnDiHS9z
l+KbVsNbKhfknPPS5ZEp3e2edEQP21JYE1MfZq957dkejDeUlr6DHVbiMyNffdYLYbViRFeHtQQA
RdmSimdfurI0WD/B0SOpjPMwO4cJBnzfGF9T6sCSuqcx/2orzvwKNJtcpnmP7U0r1NktJGtJCJ7X
4J9O5cgEYvKlVAVAnPgB9nwQ2zWj/ElARXEOswBr9AIFW6PZy9P9SwFoHtnMOKsL6ko8REr+wnLz
139c9VLup6VtuI0mUIHyY2RbOl48I+1nlHzk8iA977/+FRkvqm5WepwExBLm5wnM+bnDDbb5zci9
7heGlmueLE1fQ+xknyGquxo73xPSLKuZ2/l1uUwm78pqUbR9QjgsY19VGgruBOJ4hMJMDOOlTMv9
26N79t0cH5mv3cdW7WI5xWzv8+voV83Jd5lSvGZMSpMQMu/HumQFOuO/CUVJkz7dcagcJoVFvlzc
0FHf0ChkcxLu3yXnqeyem2ToXCoCBHsbdSBoNn54MhXY1I/j1erRQZYMSVVAcjPlD4oCah6wjokJ
hmsEgzTgQLQNrjB+zfagBkpAPWHT6amMilA9o6Hn+NcQWXXyr6djCuY9tt8XWoUcgYWCoR4MGLaL
i079UgRiXsglUYg9P74dMH1eKXcA4ukxYDJE6UUICTaNoOX/UAH5epeQ7dePaHE+lVgAZqJYlkOv
oJ/l15I1tSk/jpuOL+EfbTsPTtAu+yPE2G2b/C68cHmUd5szR71wYvIbt4z7C0TscZOmVO42vjVg
JUDTHcVXZ11oCQHAPCAr7kzVqAdi4zwwFyFSHf5rg3lWMbtIGeV2kaxsF/dcAJ6y6BHTBj+v36wQ
g/6PxZBmVGBvsfzQmL+05/hcOp1515YrCaKj6qbo7rDYQ6T572xFo5CtC/qwO2XNveg2Xe+GCY6W
rrdGCvaWKbqF6Ucfm92F1Ub511nSTNpGcVXwVO5MakCfEOaKJev1zrpkL5ilBMVbRNVM+ig/JMkK
oTkrPGAVXm0lFYi9fiOm+ac7rfq4hL92o/ksUDeP9Li6W9Dy7o4z8NxF7AJX6R7iZuRI9D2nQzRO
9+bt2Ub0RgQZFMrf95Wk1R1Kc0VmQjStwoaYUCXboAYAoD9kMr4vAdHLwSfM7eFusveUKA+E36Zr
jaYpOffLQC0xTUAUJkqX8qkol68ILnC15O5O/l29gfkf+Oak0c4zm9gUdF9RntFT2KX68IjSsYRZ
lkIDuRHYvH89M7vg0MGT0784JphUE9TNRurv5RkUnttKdbbBx95AyB/fok0tQ7ms0f3HsrYW1qKF
t1Ia5f7oZOrzcMEQB8SqKyr30XFJmI+mp7UfxHegtHlXcy7L5DC5DbqQaWIJQMHHUVhFnbt7UnDw
bZOjRcV9Jy/Qrc4D6kRdH5i3S1VWWiPJsZW1ApD4j7YbheVLTsC4L/bMHaH46NUhi0elf9Hj0Mgq
w+poxAkAdw+MatFRCt+li7h34KsLbkBbBMlVC+MxarpvMI0OXhAazjFzIAyhoNKXjg7HLzcurXYD
kGka95H4CjTLzkFRsSFCNdZB482+/F0p3ytu7FU6SapiVJsFtGlwhZjnfB2OL6lgw4tbIegcCR5S
QlsIt4wgNVKeHfHXg3h9rFBUpvzp9qsCrKLUbotz/iaGX1FKQZQ5Nm4IGqWK+sCRatmDnRZy4ELB
YpCpy1D8/cJEhtCpIrcTeHCwTJQTU/Q1tvYGqyFk+6THvUPMlX7OCfga50UGTmdxaIIe/rvzXDZs
1YsTz1ZheKT9yZ/Icbvs/M7eHcY95pMCbLefpNNGwCBs77qaC4DSi3V+WqyKe69U2sBvt9Yv6JOu
ISYUtDww7ou1C6mr9oEkjR6CRnSfGFNoK9SQrERrU7Dcd6murEcFKyhd4OyrO1TeLxcor5DrUP7i
375RmBY/+HEyiKwS49mj+XkoHTfYVY95nWbqFwEJQiFOBW0hICjLNw+9vtP8bw6eVBnPb419CktN
A5Sbt+1rIAFMFb4qP5iyF3n4uOdlVCewV1Dr4urDafu+t0vFkcjGNBIUo3GlH0yYThLRwbzqYLYf
tYVvEf32Q+MYe8E7obNlDftxCFGbWgzCFIh+lK6S5p0qECds/zpoYAtFNXX8vfgm5oPV13+xgt+2
2jxAqyqxhZRz6O+Dk5xVA9Otq1Bj8KA4yFu3AzZrqkbed4csd4dgDFwk3sHu4MTYA3GOLCFQ0AvV
1Eu0FyG4bF36ARUwmoffH2ZeejaM4UuGGPlfleUi7xbBhoglG8srn4otWhzpHDUv8YRanDWPhxY7
XZJS7IfV0M6T8ASUUSiZ+STlrBj0w0HaOWrM4z09MoodGy3T73B5/9Aq/CcBFGxg2ckTl7LPfmTb
Z/352qo489T+7o+BhVfyYt/W1cvGd7KfvVIV5nmvCfjqb1ZGkclgHfOrCrqKxt1Zc6R49vsbkA1H
5RhKO2rky55xvJj/IyN8/6LmXKeHKVT15pd9blEgOmVEAFELhJUrU+P68KnCOSpWkVlqE1aO8PD0
0U8MI6ir+leJ5Ozucjax0BVrjtxTKioBE88LKEK0+gNDUrVLTlPFBnsVEHO8CNoM5uk5W3VFNv7x
QIC0H1gDhzHvN8JiW2N8rOth5GV92LhGb2+xf3qh9tL44cCPQZap+tR/FUrXF84mD4NBPqtiFjpq
853Bavt8H1wHcTR5LUDrb8WaBk5SLYxHonPjSt1Key3jOgcaU+rtQ1yY+uNcCtfDm9QFHeewR8Ng
S/qbZkm3fc58t7PW89cdPu0j7nPmhAaDjWIPhQXg/2VrL11+beDYSvqWoVrpOwzaizcm9cPLlDZO
NliSUX7jCBl7jdbDiUOKXVoW2yRyk5YMSVso8gwYXxpMDofbi0Nn/SCgPVG/O6blD24x+TkVe3vt
ikw8pYHmBADPw/ExNKHm3rRNHM35QOKbGETcJ3FJNiIZ6EyQu2DKpiSgAIWb3Fdvt/ryqJ7QH8tj
SRTLrm54zYKsLFlh/+DePn0QHgdhlJtIM9Q1kaWdOI0RB4sCDFEaci3KCDPLucNRo19+wB3YGXZY
FpFqn1QFsfUXF47owKJRtZjZHq0VRLgGII+26tgb/RM2sSSrX0MJK6s2f8S0XcCtcf0CaXek3f8Z
HqxeufUFfThAU9bX9vWEQWVTMvklgV6aT0EMIe+K7pRIdmmlSuMIllEEY7N38MVIEfyNQVLZuD5A
mzHp0wS9hHa2NWEd9dd2segRng3Ra+NaRVCSkIcMmAZenVz7aO5SVhY6rmem0YRFkaW3nqrj2l3W
IpIQHHZZDL5CPPb039HbnIa46RVW1I3bGfOAloUiyTzLSjwwoT/ay68VT9AVeeDleVvwDizk16Sx
3Xf/EEnlYLRKtAhKOfIEywnzrxE9cOCaMM9Kmn5gdigOswjs7Zd99hIhuuUlC8qdkZxWvLD4lPq7
PasefjJusJQW5UKk3+8K48yYOneOJ4a7VQ03tsFJkUYlGLogFbm8YlpnYGIps2TNLkZ7Mf5wTbJp
1d5ex6WKqwsgR6YOb8TIZykKzhioWIQG0K847A3Rexj6tZHHD/FZk2IX3xHK7njEDO39VI5ezYMy
yo55+mX4/yBe88TWtVk26xyABxG5iCnt8syycoTxmpbHKS96L28LKxwdm68wFi8omrKCW3R3BHqW
jTkV02lM+j/GUUBivVg1nEMMJzB91QIY4M2NCqoPgO1BkLMYmIa7IZHlb3I/DA0wpBhCiPJoFkZU
tQJ4wIMrWZHd+1NDwXJG++k8iokST8O3p/unBBtVQiqLpZsv0vn3K+3F7xPgzBH1HD4zDlgN0Pnr
g7foZMk4geayYcedZBvCbhttcwKjfL4EbenHNzaEvz6/3FbWYZPkJZ1P4wmsEfpjiZUiIAR940Du
l7m32Zs0Cd4yWn1IlH6IG8p0npSzaPJPjMro4QexDtgPM7KyZxeuOrBlcWu4RfEIp0KtI9kV1otU
ybcsrFhd/KDwZrVxzdmgQf2MyATjiTFf0pvYPJ5GZXnv6zgC5DkvnxViBvd9foh4mTkV/NnxLW5W
tXY+eiMhevz73mYouHe3HzotL4Lj3wvqdWfB/qQ6/R4nqd/at0KMMbZHlchpkX1QTfqLxSyXIrZ9
DzyhXcVDSL6m3u68QNCltjeSs631JrJQh+/PjnOxkCpluF6Kc55SeHwEMHpJMxoSnP4Exi9D+PTJ
VFZhIZPdxjS5Gr8/Z4j3xdvHAW6SOOUUTFBJQdbmNXeRUCoUq+jhz3gYyTWH6/V8pSfz6dyRFJsq
EdmSHrmujqzVtBwFXjgdo8LP3bjw4pNjfoFX+d6oAVyinlx0vQOqWPXne2/78wR1/JZRt4Iz0JWj
Dxp2t7BT0E2J/LZJDET9V7/IpOtFg7Q7xwSJAXCyzB4rEH/3uoTBGcG6vq29UEyTHsGA/pCzC1sK
K1tsKb/NZOqqR3frSdAijQSsch/InsCjoi03QskRvX3YfnLflb3b6O5oQD9NieFaiQhhHOOSCyEJ
s3oM12/9VbpnNE3/L5/poRMwKxUo8hoeJ/d55p/FfNJJQgR5jemZdenpvyTX5cp+srwG6O4ur70b
MId1cj8a3hpBRutS+s6uqGE3CS9I7UP4nh3ioap6JV21dbg1vSL4wmMMb4FZmKY+L7G0KhBjM55Z
Q2gJXjKw+Au+Ct8Op/eVtpa8BkxQ89vBKJMMoMWFow+qIH3VjUpeyzNitcagg6H3GjE/tp8b1ZvF
08zOGIoxqEAvW2lQJY3v/WdCxUuPbxZDhkjUjOEDFhcEDtjA6aT/E4S1KtGbOlzR2HgHLTvYGlSx
xw0sEPIsw8UwbwwwGNqmZHPHSpUcrwhmyM+IfUtfqzPgomsmIoxEuMGrpHKThZILsL+yz2wzSAyf
bRZ1NMuF1uNWdEdbPMfhyyjUf/Fo5vIREVrER7/uBMZob6Oe1MbNSsZoc749+fYjLqhsyBCZ9aPX
RF3O0xE9JKjq4epcjW9HoTfTh5DyoLAUEy8hghTECEpUO8VftpJnMmxSEFw/5EMW4h2GjzUmCkGL
uDCnFgGDAH/oAInpgJafaDvdgDNPxzy1Ry+GoCvtl+atHJtKhMjzDg2UcaaG56vtP4Ig/3+KjVxq
h6XRlNPHR3+ZRTAVdOS9GEPg1w+FpVHXRHMFecnEqI/oIY0iEh+1mpqh76aaImO4TcvQUJjsPtC6
GRU7RA7p/fXJoFP3wjxgsK06jPz0orTWQMbLlqWhxX9ICA9E2tR6AV5djqtqwXhe2YLr6uvWtev+
2CihOfmfqxMpobYc4vs4+5lV8J+aNRNx/UC/aWn9Vmg2pyR06e63GfrP+YezfkJIsxQgXvYtUlfC
66vSPAATppUNQjPkixWt1Xa8/T3YNu+dmx9vu15owpjhb8m0PHMs9+5VA15utE9WbODKRXqtiHXA
0NwBC9MpEizEKKdUynwMKKkPOnSirYxwCsrNCgS+/rz8kPCmdIo6LZCvn91XhXQVHPdVLKCaN8QN
k5j1sYslb0pIdx7qNuNJliIV8Dbxd0PTlTP37L09tR5UO4aNZY6h3Nb0UjY4pnyhqs2QyuXM8oeJ
TX84j3oG04B34F494jyACxkcwdFdTMsoo4nxuyQU6mFbKBZS24TffrnAHkdBYe6MyuAh1dJU5r70
DWsYqsyK+zJhCmaEURwSbhVT38Q9v0OJD6QYo6v+MoGTHzP/ciaQTQl61nmXl+T6EyC8LNdQFPsK
K4nl3/CfoZ+8WCULl5qqxqY+BIl9e8rC00mNcugCi5o1dJSErQJKYss9sStZBdtA8vaEVNoiWTU8
Szd55ISGcNmkJg0x5EVeLRGo66MilkjIgRSLEo48wp1UL//Z6tQ9GvK2XgLSpLHQd6IWtAe5QLGz
XeS8gFg1z/lQEV3yFpTuxywdDtsWQIZkVHKoeDpfQPOLf52+nDlAtgodbbQpwbEKT0hlepfA16ax
QBN36joPKst6PQG8zUvf1+bHvzt0rXA087OLrTuS4FYltnbM0kCZD8NA+YgtHvzlJlZgShISe9Be
KSA3jSyYw2WQrqFWjOf+svswYCgc4JNrwG4wq0TkOasEKFsNVi/x0h+RsIlzckaOW2ncZC7sDR3L
BeQjA/iG5qCu051fg3dMKjVKqgHuRED29D6C50pVeH6ku4rJX3Uc02zOLuvlrCnPO1AW35e04e5s
XTqJdqnfJFDt/5VsSX1Zqm9FUCw7hlkOBsOiV1cGGmdwk+5mUA5dw3apmq9MFbu8yZ5VxfK5l5JB
MPie8FWW+pBJyOs5FsQDQvCktZzQerExHGHwhlhHn95k5PaK/WTfGJq3UU5ZeJQYTsFsXZ2mpEoV
p3xYQxR7NqEbAl7y94x451/MtRCsvpfj5T0M7T23FyKNgH1M9O07ycrulmCO7kcKh6l+B33Jsiz6
Er6YmweJD510mr9NYJGqaUh1scfuUz4PrP6stoCYj9rJ6nIEcoG4tjgRFchqpi+vq7vSS6Vte7Hg
8fY4WItAAOLsK0NtyetS+jYb4q78XbElRtuJeo+Q7zVXfOTQvp79YF3Za2SnGpUYj/pG9a2N7VTE
3VKFu48a/j8djy7LpgQc08QAYUygz83mqG3KHtNnG3oEgywBXTv0vsamYvZyk4xlpd/NAIKMTSSE
wF4Y/YoPrTZiAeSmeht+uTVLj+lsX2oFt386bqsih2hfKAnaLhNWt5G4QD5JFOpCu3n44wisM+dZ
ubyfApXY8+yDiID7j13jTdbgwV8nps3ZIlpaPXMpfsN4Fgjb8Wdc8h+zbUn7YKNxiEBxCoKJZWXb
Noh4zjMr2XUX40Tdj+IW1yThgM4ZAYKWm4P5uVo/QDjLhPN6S9xoxZSru035Rn0Lph+jTxsFVeF0
163yWPd819e5gPgzU2l00MSEOE+gBVpjv6aikmAouIuNWjByaW2LR5CdVWGrhv9QFW+T37oBNGxT
tdTCu/DKHO/mT4OZaKI6sLGKGd5f+uMIPkYtc8cvBN7OzNTYKhrR85SeDO5bfeTjQIqGyeJGGLsp
kOpwuFBbAgwOuXwitz6XRMru/RGqw0ygJdqLU8+azQkjVEwC94PbWQPdmx308v+Qmhl8otM7PL1m
oVm5qJpe/n+D3luoZDocakHMIj3y44MkUUaJNNxjoJhnaNaDUGYv+7iye1MJ5DE42mAiZJIyIIUa
8+4MuRPPk4q5ruu0FTarO0w9GT0OERWG0tY6y99SRnrMliEumry2pbRU2pYng3STegKBNQTdFnnr
9OYxPK07Y8KGpyfGqPOkVRBMrt4tRIBvwSlWA/2J/bpGakri4WGN28zXpnGX2fX5Ks9Eiow0GQwE
ASmlnCUdTNZHepyj9hhbUirbZoVzE5FcPPGMZTpnWHAkcavC9LaXDfFkICU2cufvbudEFXcriXGw
1wYjzrVfOQdI49Yr6ypNHMet/6wP8RKDZ9856LJ4qziDt7RkNUM1J0ocCDedUfUaV4kECQUPn5g8
dQlBbwSZ+7Bwe14fgz70KEZjDpFMXYet7qtCcGJXBu63V4yYHQ64cmSfZeDf2j/AskYTvR75KpIo
CcePrmT8kYEKZTl7PTscgPIraDoQU62k50UvsU4oLC1Wn0zAFvZ7vlGfMUjKe0Db0rNOt3hCZU7M
A+trGqZp9YPs5OnEeFaK/xK4BK5sQvtMIbLwgPOmFynTbb/5E4wGLON82xNoJfSVDEIdhCbVT5Ow
ysTWXBWO9J67VzKcUqs/XTkD1MF4Zsw180RTaQIm8v6AmQ1mH3C4JMS/u4anAVGPpms6vo3XlgZu
MQSyl356zJGA1owr6MJpTKgR9b67rNmkbtxp6tT6Kt375uQ5cwc5ilxwSNz8TuAopZi5FURhUco3
zoQClC60hGWQjcEINBaMYbkzX6lwc5a6Z31xsYabZPiXu+Biz7NYpN0VPRo6MUn7CdqNyfXrHbNB
7kp/Kd5EKOa0GsBPsiFdB8bPI+HwVoz3vq7prt0YNd4xiwRI1G/fLaIaUtnjtI9+l2n3b3NkR3Cd
uNGQ74HVbeQoDC8kiWRgWzyB6l/LFMS3GasC9ZadLxBn5ZcyQzMs1gi8dPqyLDIAsM2uj88WsgGy
R0VLmqDWZDfjB/8JtRaGcjAI96trWDyNkMtRctGlvQp+bVJSI/JUtDasaHfNOsdImGoZW1wktPYJ
hMJ9qUrtK6K+N5PPL60W7gMMj+x97aWo88k8UXUnOQMgadlsS/GOWULyM9II5X08Zej6PUNiYSDt
27XkTM0ltw5CBDpSQm1spNNXCL172gQgNVWW9VfiNxYuNNfCzYLidsqT++BBuuEvKKrHIp/EEHUK
BvG66hA/IiCRrSFAGwaulDPVqR7T6uelLhoR41uWiBxftuxFx6O6mSi+svPkGiTzmrqUK1jFfEoy
IVPrTFI7FzVjYL9RLw/c1EIOLGk0pDAQCgKtujbVL0f9Xn9Dj0NDdYOU3edFgFbRpGsjoowDbeTS
i127I4f5v7fOGO+csWRBzQLDxfpNMjnqqUc4HkKiLj1kQ1m5y4Maz7RouYaFiiq0gbwwXqh4TKi7
U+PYW1B61Eo+FAdB0Zp2bYfYazVe/H870uuKexTHhcKflafAMwhbPBvmVLo6aGoa67xD8v+xiHv3
Y7aiqGu0AMBZKHkqFS3N46WvaFOy6IIMZZWOHJxuEdpcCC0naNGYP4/uQAw54G9wipwQt3bBUxav
V/LhVRPmSm2qKYkrPYvaoO9mO/angUDsbKau+Jb7qQEmGu7k0rmpYajWyvnDDpB7JEHKJIuBcRh3
FlmIm2eZGaYaR2W/soG4RZiRDNyMYPE9becKGJN7HitllkMzxx/t9w2GYNhou1NYY0YbmJZqoyp4
9fUlcG8UYVmkyctyFsDcn71NUj7D/WzD5JdwkSfHR7xaXETmJV/uTtOd2sLhVfZaLQpQg75Art8S
eXugxcmZkVWVloLDXwHDfwaH5gABAHJh3JmpFLA5LAJB6JVjS/SKaF79maPTfMyA1iiSGIwsjVrT
kwCqYg0hOPQEeqcRFYX6LGqY2nAiAsQH39Ja74R3l/abVmA4+DmvtEKKzReJ5zYYj0RDrZ+nVI4F
jLL19CZJJQ4hCc2DgPGtbyEH3qbJU2deZswrTNi2yNJN3RLz3SuTkoM7oKrdEUjMviYl5y19UGEc
LDU0hVmiSYr6bB2RyUJzLyWsXCY5A6QsPPjVp+08FKcd7acu1ca6PoPEQOS+tuHOIM13evq6L8x9
n3l0QW9LORnI7CgdcUDj9nC8EkZX3gyU+zJ54tTmKvLph6vVcv8GVyKiX0aPpp6woBOnlTNZQwQj
dO8oN+p/2GdZw+/SZmDkNFnUN0EfsQZWa7fHoaw0myQUMlKPnivA+qsPUcgm9WvtFVcVy9AjnRzW
GSa7w09mdRrOwB5s219U95/UKDIsfA8cmdT16RDFspnJW0jmLZ48z/y46kxSB3SlhGiOFGyu28ve
jaQdiPPhAjVAxuSYPIXkmKR/leTU5EVdtjgohh4FEu3U3ZGnhXsYVIYbADqvA/rSSTXhxVPn7jyj
wEoA/3bruugGng5MHYTLMu3e023imzUQHgDFWdTExfhaw9nYyrT3HZ61YMcobPyJ3b6Edsrldw+z
VwmcdzBD7j138eaUv12rNi1GNL3RnfmS8VKw2nKfF6mICqUPMUkcD59vFhi0jkJlB2OFHtRhGLOQ
zIXo6susLgB/lkIOC1QvBUo5O0kMnabGb3zCRqrVbM8PL+QRJy0Rp9e79S2RKKKMgD6z33hEte4f
BryBmcZxydPjHilUTSXCcYz3OgK3ZJuKiUg8pzDUzmElazKyyi3seG309RZSBIKOFgir4oSssPEg
yOo8ICRXShQiRZJowIekTnPMNxRrfQAMYmVqTe3jh96oakYRsNsWDBmcOOI4BJpLyqNdtCpAxN+s
5u8OA++EVfC5jWQtGHjC6m1F2sK/l/hzlbFkPHSz1T9M8iaruulDim8J+Mi4TQPKR3wpKN1/ekrW
7v7R7rNjdYN+fWmR/1gi2S7e+z6d4g1MZbi9GxBwyucgkTA0YvavF/NzsDG30OR7/zEgoFGlfyXN
cJpBy6WYlTLI3wt7DjFM9zNV5FaTPR45OvH0FHWph4AlHfbbB7qG52oZtqVUD29phLM/0AciNGCA
fANhtt/igSzTCBtq+kFBShUf4e0aqfiBLKfrCBGrc5u7lw96xNWaIihbSgZnQZeAPzuRRXGl1x0D
EC+u1qT+V4vfnFuPYxhd2pBG34ce4nK5KTuNpHQaeEQF0qJBx0g3GuN/RXByI7lULFoT4GNU7dNB
DucuEMI8i6T7keuJhSP9uzbAFgGZmOLmgwiGkCtbujo+UNJITYX4AzKpGesIs5vfWX4475mTbKCx
uDt174SIX25v68b9NIBAyNO7hDuhiG74YT0jaKi3H9G6xbqXroj04WaAkZI+msPLIYoqj1F7XiSd
uW246A1qyyL85IvmhujwWgLJQYDBRBiayM9F10LinMn/o2yyFdv82o2xg1bx/0k+Z1ra4Zs1v1BB
+fZP1JLaTaNVdLJg/vlx7VbkvMEOuy3x+K/6MmPWlzNZNLztdJNqAu0+DHXSYNE7io/rnCmeYQAm
d9W7/5go6uAppmT/IVL8mUVMVpC5EWLuo1YdyYQvijY+/O8KBF6xcBmgrBO6DdyjTNyAkuuDL33b
e8T/P3GCZHJ+7yZEt9EAmo/g1GkbpU2/M0X/uFbIS7bIcX1CyyzQqCwXhc2fk2lC88bEZjAzYiGd
XD3L0wsATQDQ+do3YI5/nUKRYE+I+Y6Xv1RuOmsNCMGm4GokGQxNHVk6Nm027lKtfUr1DEYIIZSZ
meHKrQ8ZQU1lojCn+bSbuXqamvLiy5a17ObI77Rb09YdPpYVm2CjVLF1Ra+qiSvlUuH2iqO10kUD
o+SezpvrbJyByMWnGM+UXf8YWHtQ2zC3m61pogAEXRK56q5GCKX7bQxsT652aOAjR85G4HbfSmF7
UparHPDpkbanK7mHvnHrWNuzxCBxr1FWe2mA9kdzBb3JI8+mQD4wi2+/NAAC6ugwYJf9Tf7Erxqz
rFUpkYJyIUyuOXsKrXQW9QE1esei05ol5ecE0GoBUne7biW6muZSOd5EuBf1Aon6CxCbRiBJU6qz
UIfeN9NNggK1cCM6BBvI/qu49RhhcY0/OJVUKTDFhjErYmUkieSJyeJleHsrvt7yD0xZ0LoQgdI1
fJFTHgqDTYYzNxYAz+TI88c5SDivKcQRnJwAqZelmZ4ljWmp+x3jsfOhuNfxJZ2IRYii3FudA0Nj
uu7/VtU94Q1reeh9QNmFfOIbPoXK9fTmV5RcPnRuZq9/CySY7xP/gB4dxhxavt4En/kj7Y4mdZDE
6S/tZ4IG3Y7rHSeNrDuo7Zk+caGXRjYPvFdoPtOJup/H8XlHa0orMq9lqqk5sKoEHQNWR1pf/sx9
NBdhaRUNkTxGMJjgdEUqhDTs0ncJ1OckswrjuxWd6Tg/j1BhLVdzWzdaMjMWiLXHpwouVR2nB5iq
s5QuSWHGCTPeCE4RK795u6TnaU7b6xd18RnfLIKjSqFeKkmm9Ju5teGGdhe7NO6VHcMmILgsE3yn
Xn0VuYn44FBjw/d8KFyNWmcdfv5D6S6XJH/72wJuOsx1enA7TfYwO4wGeoqLSZL2ybodjjPbU2wr
waFyIyy99sa4hQRyT5ews5k3dgpzoROTycS8wDqHmZMhESTPNbiDUXumwCYm9pKkemNlSBoRM2sc
qCj3WorNgM7DWmikZPijiuapFb7J+fNXTgRa8HXyyo1HWX8FTMXcvjW/wcknELrl2GKKRMiU1Ojr
zQT/UbdXbC/T89DlG/VJQ9Da9inJOvinm0FlL07/lqI0zuth+jmhoK46wTfcIgzEWnzV0WgCgixd
Q3Scf0doy3QVAqB48YCCFAfffNhpgUIPApPemuEYNRQwCDDi6TkZYbFma58YFMCO1hdR3SMujoaU
monZIo7iPGhNv+T6h3QVnkfiaBo6h+7S4z+HmqXFbp9jrcrhZwT24VCCVo/r6ngO1NCtrlRwgLhR
kWHf5zxv/8SY6RUnUwmwVH2CAFbD6QpKEFo6+FzxoP8a3dJqIbspCJyiL1BppMg8Qdn9pkpQUB7Z
s4W6vslQmIIsY1GnO3DHK9EKV0E3I90tSnx2vQFhOr5vh/BxiczFBeLav8p+gspgG4rRrpJI6ZbI
FWv51MOy+Xexuss+RkL06YscVFXzba16LKSMgdIoyIbJKS+y64IKpmD6jp98n/esMuGHJhKl9KJw
drsL+3wFc8lj27ZeEdC7qYUfGsos5aZY0HmC0YwF5mpHD/QvuuC23zOBr3wosBsTQpB8fx9VuJti
HzPIthwsapwqI+FkIENfxrakDAAcW5cYFA+SVypMN8EgNMZs/vLZUtR+N04bLEs9Dl1d/9gw0PMA
gGyd5e0wnJL3MR8ln6IW2ySoVg3ZZTYZHzo8174k5kIvBc0n2I5iVWo2cfe1rv6s+1enOLiTKb6U
fC6AWdMPmaP+eU1N7Zf3E0T36+qbqRK0c8J2uKFTDNr5L2H677FQm4rC8riiYyKLlzcrQRaHAO9d
O+Pyxf9ORGn43PwNzajDNvfdOyFyTFUZTZm52jhGm1z5Sy+zC33NoZAt7T5Ky1n2SWIXxrcZXKdQ
4uLn+c/s/wHcvV1YaMHVHAf3tRVh8fQaV9iPXtlugAoJworbYXQtrd26++J2xmPZMV8w8Uqdra3m
gk2tdCB153fWnczqB8ItTufahYk5C4ZCu2i/VrMLKrEPXMmXuJDsZB1qaIIOCOl9sJuQWFndi3pF
oUmN/FylnEQFJFY/G7CCLWKS/E3AQ0LQAuuKOZLa80TfFWmGk0UTGnuLWbgFraVTFm1Am/w+odj6
F2iY1DnVR3FEGIHBUwn+TiGTZuqX9ij4NelI9scBSKiM9ZmbZKFmgMRsNm3AYyPxdYd1LkRt3n3I
NJFd6kB+C5eHnhI7nzcSICbKPs7w7aXFKZXVkP662qRnvPoKZrmaJHKikmPb64Bg5TpZCydM6slp
+IxopdxUPx7H9AWoUbUZeCe0NpPBmWm3Do5eiLbQ62M1HjppHj7MLbLXcvxwF7KI/fU3kPxGxSJ9
nENtAb7Vgd1qoeyhYxHsj5edU+sB0imgDWECSNHe8luOjMhglb0AfQ/L79jTyWcYDF+Idlmw47mK
9u3B0aTtd9YmD6xRaPxajWOMqYOXmERsCzmDavzOwhvOb6eNO3rXI79mkMc4pOnLpb1CP4F6gKZm
VKEqo1Mx/wdrYKTq7xa9W6+mU5+7c2JKC45StZfx+XbiORn+14L9eJj0oCEJ0r4cDBfQADXvdWtV
+VN3dKTOdS5uZaFfL27ZAAY3v2sosufB6OM2cTC96HtvU5xLPJV5E50rqRu6J4WhopzMy1pnFVXj
ClwXpwEkeSvhZrAWYAIUq3CdUN43RcJUfz0sm/fx0kpEFMtrVENCgBeTUb2up+YubDZAfYhGKTWu
DM2ZZvTpdkkoWyksZMlz+LFlncyEvBSwc63poi3aLbc/hnTIFJwAKo0OmXjagcGW7bydCkWPlhPI
+2q4BEkvI5/jmdJ7AYdWwGApkBV3z6dfIsTEvjJ7ciK27DvzQUyBeMzwdAIN+wtkjzXyLUIUuBzK
d8TVeo0cc45g3h+TWbTy75X2qM8Ize7yu3O5qwHoipJgCfVcXH2acUfog646kdnwtzCQ1FRHFDfZ
1u7uzwgZRDy74PntFJrIq4p5W8Ax8YqoMMEWTXPn9LbGn/4/rHkdmyQPNP2yDahegl6Uxr3UsIi7
mZoADcO70whVHzh98z1y4flndJxJbfd4/GRL1PKVfA1y/DHghCPtMA/RKnHDBiQGUgDhM9xP81nx
RWkbeivwZtDjy9pU+bEGEfAcuayre/Bx4IQyxTgkCOYcrFcX3jCeyurDlEGCoOXFVCSGkqhvZ9lg
5Sh1SCjNrjv3CnhcCbx038fch/JYPrYUpSt9NJGBNiVV4ffQD/KMOSsumIm+zUesqd3iXNu3TZkY
V7iZu78PhEb65gEEm7d0M+M9OWj1qRO4gB3d+YNY5TTNDd57QqybijI4u0Jzd+xt/9aNSjCnE3oc
sP6Be3dEwXsJWlzMizxi2Z1uezE0ldIUxqR3uAjEmEfBN2tKZ+P12qkA+5KhzYIWWeZTy7B+/kRZ
sd2anRXiNkP+8upYwWskpujoXPN/NoZ6x5+HYfgB7sOUzMIT5oPEgAxJgrLciq6CIKm0C5cdXzyk
pbk14SfF+ZORICCN+eY4e9Av+ISYnb5+2V/yM2ZuugE9/FZ6L07GzBQU3g2+JbD0ZvRI47Xbowtz
UpR2UiBEjlmQTJCmHCqRshP+H6r21GjHGAg/+Xnqh/NHOAkKZGNrc8v1UMIe8FxCAXNSMheFT4Qx
2+onrdsZY81bLu+8u7XrUNYXps2jG1WXSrmA19isGnVBEj0fzko6jrkJHXiGB0otIngcykLZBImV
gt+9G0sut1HxCKM77kS+HyEDATJQlzS5hNoswlSVVzYkepB/x8ux4At42GPbRvtsU0Jc0EC/RCVC
i0BY/EdxBdy4CRigFbH6Z/gThFxLzuAJiv/wUHkewXMt8XypSqXDytFRtKUBKqu9dwnGu7JMFIrD
mEScK0D33ecHwNfBPdV/wQiFlKJBfXKl20P37wHKVzCd178TGGE7I2BTRsWgKpVy2JQkfnMxxFqV
8zYCrDRb0JvhzlC4+d1CkUOJRLIrI6zSfcruBavo7u2u3vrcmxta2WiTaqRmdOGeDgJkj4kCZ0vy
wiCJ8d2ZGevk3S5NcpVEwMq6L6NbJNKLxdIvrUJl1beJM3t7NAVrXYImiPHigNHAH8P9VsDREkNX
axAepRTdhOmEJt46H9zYRbVumAOPEQLlAGoWrDPBs84IevSILsmdv+ys81bDXMsa/JSp7EvOH8G/
1L3eoi+y/F1JI33euU7jcfKqmaOEXO+srGVTxjmKrk/GLe8OJDVtyMTFC5jxTTYXG81CrPTqof4T
aYGqjC7/KGt8t4o/59q2mvr1vJ1SvQs5hnvFcSnn2e6VaOAZseCBKn72nNxsPIEaC66dwUOP/69g
Np9pVc9lbT2forX9bCteov2HXzuArDdWMf4DYNYS3jwW4qDycavPVjwXNGTUj1YV4pUgcactE02t
84pUhZF4XeH5gvHwCFJabeY+zcEIXPXl9qTjOPhNJ8h2sGMu/RtUZtyOI+8gXceKNlBNTlyfgDoI
pnkW2E/UEbvZLRdAfl8lg5ic0rGOCFzkTDEaXPfCacEelxMTUEIEy+iq4ms9EGyQuRMjeqD+Rq2C
pYuw+ltrpdHdGGnZx6l9beX/fvQA2OuYNj+YYVBp+EN7Zgmkb3QebWTyX1DJZjako+mpbOSxzIhE
2iNKJ+agaV9A4PLGjrN/wZgdZjzfJ6BJIZIO4Hb/illUDVm/A7NlxgWMFjRVz0n2CiWRoopDBTIs
HUDQSJ2uOlr9ahTMlsYj3HR4uG5hlB47hPcLXW04FuSP91YpKveL1I5w8CRKthyu5ToDkWP4RTQ1
VsTgnFBrsnEi84Acn8Kj7ay99fHIBuHVSWLCIBPGeL+KP9KHocZLP92KxLi68mv/fnCdgA492hjd
QncOmPYeCbXmdN93lizODvfo8kwk5f3UlfclgwSxkE1DO7jqaJ8a77hCpExFbcP8sHw0XkSVxgGe
clURDPC6k8mQCVYVKKd6YDwQJ9x5yrxEGl7qwXv/KT+wx+IqVgfi1+ToxDMw+BnGL6YW/xnfvgV5
QnuZQsMUeAYE2kVFincGBfNRmNUpTZKy14IoFCfSRpRzMwvZvXKL51jha0ksPhAdP4UpfwOoI6l6
PintrDZrccbxfgVIi/yqYL5djskV44IsbPDXlFqiJgH4loS0iFUptzOsRTYoO/jkQZPyrbVi6aaH
Iu95Io8/0JAmph2/a248Z97FZuQkA0Ylr8CS/db6N3NSrKT7lbG9ASiTni7RzvXr4xEQ/iYUXgEo
9Tju3Pvr7w9XJAj5KcnvuWA+l6EqRdNzpLhpf7zBELJobjpkO/cyYDSBvQxZNVdpUcCSERyb7uYB
i1uMXqhqT/2emSJo1PJMPyxLa40pqWgIYvJovc4suuu0oJK6ubYc4zW5nOSaCMNtS6O/BxGRODup
77lwQ/AtVu6JCPOpimZh82cAAl8zkWfEltMb5CMb15dVcoMeizML2HAAYE/QonU5bALP1fAeCsXM
DfrY/JWJGqWXQuq2UXxT5dWdwm7dOiCk0FiZEYgaWg8ZbmL7zXJ2qWmWpD8citZWi0nASr4xGdmN
lUaF1/j34buM0Q576wg3Ic/rItp3kzxekcg20oig+PI7JpntO4Tc94l6cik5oWRgVKaE5jHBJQAZ
HPegj7kj602jIRzWXvbab9OAwPTHKT4mT3xIpqBtrw548ls4w8muAiawZoADciJ6UdrVa5ev2HoI
W6D81z7qF5CcQmO65ITXXuQeL7qGM9Gt462ha6pjFviY6xbLcSb4zrSzPAcpMOCjz6wUPRkwfMNB
8389SScFs1ju4IXhE4ILwgkPPPlmzwGtGjprAjOCeHvyUvzFp5wgMuida+JBeLlAZ+iGx3Xhcdit
22olH4hf6x6TqwCB2iaOb74PG8e7CPFbXiKa9cXehaE6wtNeqAzKwKatO8o6GW+b8HoGHBFlBtvx
XSBi4IIbYHYoWhIKQpGj4diHDHszPb26rh4l4SakFMFourwGk6UQUhBXKezB3GhhuaIwsLxsUcCU
bcprA9IoTRJpv9BttZYI/nxso7zXY0orSOlZcbtE9S1cPqkVSJBl5WTev4/sZcQdsFsFxfZT+Jec
8nIVU9S/tiQFH0YesfQdkhRhfTpaseWidjOKytC3ZpUDTTxzOl9ouAps18hOU6656yF4vsSTbqSv
+yLx3wCUCzBfhhAATULRSg961S5kwCPxTpvSgTCOR17x+eM7DKfWIBvH3bAg2AsYysEjYz3qOQAF
rePeVhnsaAidk16grwT4Ujz1uj8SpYCXS1pVGh3yOv3QhxuMaFA134n2MZx8DP6uS3HmwGScNs3b
6+9cDcnxwENbDdpetzrhi+rNh2ZhFFD1E/rebwPLvhHf0Myndt2EFbU6PBScDsqgT51FS8nMTC1Q
FA4rlaqqkfNlkNdGj+tGOyGRLqBDtOz7YYRX0y8ivsMr0mP7WM97I77zQET/UZiAl40aUcDpEUIS
D+Gqnp+pouzXy+X5kKDl3jFV3h4vCuRxIrwVhmnOQCwicIxzLyO6V22cbkGxUES7U8+R4JDGyuiE
oRc+kcZHAKw5jJS0fZktEagCjpOzet3hi6L9XaoCORrpV/NQZP2T7LYzlhcxbwmADH75EjP22L0W
euAbTZCpCogJnkmPjEBopbWEPUv48SdJv/Y/iwVaH0MaVFqpCp5g4pVHS4FFo85FBh9P2xY+9V/m
0YZlOaPlsccZnjXImK3MRcnlu0hdkfz2qANlM4mnUqhUVPSPyuSqiarnkqy6vAlk0eSdAmWwMy4K
bf0wTj7hTyJhFLdO6B22oe/X8xqibWMToNYk6ap/KcnQBiFH3+eN44j51hBsMjevWSn1itFiE7Wr
ucRuOObTQqQLMTvpxVqMtKeIqZM9UIL5QIY8+W2yTkIeLmZHXP9ACQXpo+SV8RswpcMaDqmPwodc
YQ52dFp8aPufzCTkru5xmvZ0jbg36zNULm9+sIOH6vkSn1d6A0P2MZNv/u7+i//e0pbsoCknOtJ0
oZ6SUGMUnert5I6ASDLD5ekHVNSCryPbV3H0Euw0TEGnlmkf8kMH9Igo1mDCa5E8t+IEDKkVpaSF
o0UN/afPq72ehZLL1rYkEN28OTIJGAzk55fzEyM9E+NnV9rPVVj03ZdSNAobM0zq0FFYUui5jVUM
VcxVR7U9LzpGXUwa2gKWCkXP0kR5i8roTqEg5XJ4aeg/fFk1T3f7CL6hXTOdBPnX/EBCojad4EJ0
IEVWFowayDwHlkuAXzlE+Dj8qU5X5sQR980D9ZZz+kA1ZlC+fxoRUbjLmVMyZlvhvdhSaDRa87YP
K3lpEfUcGoZQPs1mLqGYBj9369TsGtzBU6PVkQwCRZDTgFNIYSugNjx/77VrxPHGwoaKKgB8Q3bx
Gqy1KIJAR/CUKdpKr6HTt8vyP6qyOPM9AFvJXNWAAqoKWAzeaaFyONFJpHUCaTI7S/DmvknEDpwm
GKfVnQ3Lf9ffDcbIso/IVLCDdoycOLS09xflssIqN/+/HBBzBqWPa50pUDZ/382QQtxL2d2o6VBe
v5PcNk18P0n0zujhs9nvQSrqGmdZUuq4OoBDnn2NfdBIHAOy16cBFTdVfRXVhZ9kz9g0u9uiPF+i
IdCnFUEV2GWN+wXiAlrBj8dCJzFhQWiXO2EMr+ZebwusSC5IF6FD0YuYnf5bcAknr0sVuUpftHcn
llyR5IyUl4ql48SuP1jerKawyg9mrrkQTJkm5nl6rhFbiPPBYRnGJomXNty6qucAfrPVHeM3mWEq
nKJApHLrH2LgZzcX8AMfEa/xNzM5iA1XqLHk5W1BbQnAB+/T0QiqTpC41wodB1VVrUo5ig+p/mnw
no62QO11QTknoND/hBteHmnwRj8kCABDsO6c9pj6W2SGlpN1YjQ9qIHl78bAARu/DLdKB4gyNi0l
ZwgTqQfpq/J/ES8/x/h29rsvsow1E/QV4phKAv0+LVa8I2v18EHD6uULuRIyWoqhMWpYrkMYcCjf
tT9srg11H10Q0FZpKBtnlr15qlJLItAUoDbqZnpmA/DzXAok5Rnv7zR4a5Mi1QlMxJu4SbBVkjLe
/r7aus9mDYX4s4sKy2LozkUq82WPYvQ+wxoffyqHvBGv3Q8RoAK1LM1n2ziitesE/mj+qwxOyrZ2
4z5Br0SkLFRNpnPYwTBjmuERaDx4VeTvFl/LlZoq/cOT0i9Fajc4HunS1yJoyE73j5fxhRA0GxqE
4d4FJczaWNIw2PCxs7WxTmdJjB5sI8Tj7UoTVoyqFoJAO24OGAfKStHP5fOqSLRJYXQ7R5+GbUbb
BNQsJ/Pz7IlWSIPqw6KnbVb9FW4mKxayXfjmTgPp+a4ZSjuhgnP5EsspllTjOQlL56tPiJOjVeR0
TdiY7/UezozJgCnyttXlUBypm41Rub1UZmwcrijlALvLCiSXjHEf+HSGIHAlB4vW6MEERlNDg6J8
ycFC3iTcxMr6v1ftmoWMVBXRfX77cSxz7dCVUVhvRFpjAWA2AEwCXtZXMVMkhtpXyS+n/wblVwD1
9zb8ArWLs/76vBY0FzrrhFpledkw53D538a/To+bhnijHQ1rzDOdvOxWyOZzwXb+6Hq1Qm8QkIZp
w7p0qsoxYKRjOpNiHVgOkurN8LiRfAnNP+b5TCPZyTuSHf34bXZfEv8EH7ock0ImWkTlSC2AjJ5b
KrOiKoObYR+t3Qhrp9QPeNRl2p+fb2xZhKaWh55UgsJDow3Wx65B5dEXVhoGwh05bB4wQLL8WZWa
3rx7ijeMKTjZoI8Y7Bnh83tD141PzAB8ag1mZXBPldL8IE4zaSCL0LuJYU+F7R+cnbxdxXQvi1k5
ex7VV6hiI6N0S4WB85O+LIaKJ+UOQlc0PL02HyCp3lG+PlXrNI6c819LQK0c1XBV32u55cZLFt+o
7YHSOtGbgFIXRvRI0GasIrwpjHe+Zo4yP/J8ixCixnMhx0ZeaEx3bWwGdL14auul5Qt2W7WiSJKQ
zJdI3hXSH/bJHyQmjhv/zXOlzr0Er4QyDz/JXah7sbu/8mN5EJLq7nf05m0+cXBAHp8Ta6I+prqA
+kUK6PIasI/1BTaXFiyBjt/pVIk2krVB9KdRkSh/KQgdHpfGvwgRbj2kH2VzIFKr2DjfNk5eQx5i
JXW7M3LqQ2AnMPMfeZf2ltnP5qiZBlp6YKPsTf0qsA8wexeIc5E3ajO269xR62zUl5hF2OknRmsN
qhVAlqLo8245GUlpXNkBfWD4FV5cNQGNDE7AJwwk+PK6Zj9XNA8nQ6RfrQPgPNUQpoHjq7fbWa04
zbj3umA4luw5983Jr5YTSR9WU3WdZOGwYRZS3c/lpDcrV3gQuOpQ7gHK4JJs5RM9wCZ7NFNXnTmv
UKASq7Vua1myr0iVSn2Sc37WwdCtkzS9eY2O62HyePbvqhrtm5p7QuCL6VGd69oOY1OhlQEXc1RT
dexwiMXjlIlIoroQeWqFaDSEk/RoL3WMVEr3QQaXu1OiYuw+9qHh5K7zfbSOmHXo9n9u17UhpoRI
XD+fKWUQhznmQ53oRm39gQLpQskIU0/nlCF8KrwsZgal3IV+XC2RVlCuJBJYbHRJvf11umFiTSkX
hJuFtU7bAWPiJ2kdxJC2ksaCQMS1Q+w5LQn7KVTuMM70zc5RZXf46PR38BxRcmlMcMNyCA2rwuyX
ucF0GOXoftCK4bm92i3Bi/bg0NwwyJtwcQrUyZNcyubUL9IvzJWzmoi3Pj5BUgiA9UC9psyCio9i
7KK+spMefCmSOoJQ3rqX9r050AQnhNial09aB5m2zMSO3VQ3e9+t6m91igWMzssHNz+SW4UpP88K
CbPZLVu99gTjPY8sg4s9GObyX+mdZK0NKZNo9dA+jKjWPc7XzgBsLPa7bkKBOHLR4puIITQbwc73
rWAIFogPSBu62JdbeJZMAAX0FvDjgltqJiV5oK6L/mEGH8Bdi67iNpjDxWE9KywGrAdWZNI+WxaD
PdFwTjMesaQfX9JxBBpAJ+h6oXI1iDVXcRGDpLy9kk3XKU2cMNEbLNgLlKywoL9xzWNihRWTHITD
PwXsOb/UDFZKvBIab/b3QZTzIM1/e1y2HWRJJG8eyQUN83rP9XEhfNfHAguaUWQAtPgdGFxIMgJx
/yQPf90cWaaCkkfrtvIxFVVmATNFYZHskKkAN/1NuPRQPgkJRY/sh1RYHelgM9OdcR6uh/OF2QK5
FP/Onj6j9IelT+mrG7ZX39+tl8cBSJvS2QOsEJSq9zAtbDDuOcBoLVih1iNCwzhZdNJU6BAGdNSa
/C5K2/NxlXwQcHHCtP4DruLlHfoax1coyQWwtkofwbR33Jm+cy3JtULTOVRCdtuk00StdvashMBf
91HJAWe1wEqJUwmW3ZtKeLUqCshcqiL9+sKesEpip6gTM8K037cxun2v1Hl/oGjkRuF5I2a7Je9q
LNGkqYQxPgnEWcF0bXCjJzWAQRCcNwb1mRIG6A9Fxcfniq/BA+ZMIiISw/S3cgjAdEoa22E9Qi+q
GRo320fr0V03Sq3gYK8/znNqUYGyYdg7lTXwt3GXRQAumivXIkfZqpKwTuB/AzL8A7djxTdVqMzm
8Fv5TzMjgcXSXpkT/AoVLbtZRiGo34lUf1M6zxLWkyXDNloA0e0oSpSCcBt1h25WV8zCZ+B2Bcbt
EHCe3hJYa85q/PzsDLXniLGR6KZP07/8ZjNvRaaLrQNBwmgGCLIykIfANTR+dV6BL8h83xQeYMwa
6GM5qxASS2c20jqGDUwcqGsuh9NBd6fLKU0H7f04w9jrOBHey2u0VyJ50ieFyC2bX2U5z6dveNQK
ApfEE9RUy4QHTnwVwEoduy5Pnc6rx0w4jmL5mJtuJrol5J7fLzbN4+V3fAcMgo4+h5ZNBkes0Zme
a1UuI8F7NU0a1y2eWNhOctaK9b0/lWkM8MMC8fAcjGr2mN7F8RwJ+GRktuxHnOwAtV7KldkFor3a
Ns6JKIStLjGXwKWzbHCy8gGGOxVm73AcjPRntKx9GUMp5ikwHlzpgHSsTY69zLgfQEf6okjHshXN
EEOpx5v1JoJEgaHmL1EAY8uXnz48xyXCTAwI2SKBdXsUAct/B+Hvh4J787PkSr+od7wFSak4LwFY
DjuKkkkZgShAq13yJn3JlJnNK9Ak2GpCZoqHUkCFnZP6A1Kll481pzGZO+gx+Vxs7vx6JjlZOO+v
sa6Lp/dxm2F7wvFMfEmqbRz0bH4d7DDQFx5zxnVK+SpTHxSieeaXPg59C5x17l9u2wID75jWNDdW
oOD4HKTOXb+qEtPBTUBKTySqFE+MTGLyrIhkGtcAAWVWIMs2vvHbwjyrfvHz3KWj5MMjKx473DpZ
RDUg62MQZRamNrMmH/9FODUiRBt4JWHqr7/HO9xc/t87EtqdwtJz5/2bx7rVnYCdoo6xwQHXAedk
vutRTsfX2FnzbOUiNCAuzJEMY/dtdBZ/b9BSOFHmC1ThPYxRiADACdTtNjKGce1Ft21UVyArjP8Q
lUPd5/YYLaqapBdo91A0c90X0ocGCFuz91Jbkmx6nLHoQEAoQSrCR0+eidenPG39IiO+3s+6g3EE
dx5Xx1FR0Ozqyg5F1/8CqKw2+EtbFJDJbMTZecs6rvKihliTq1RmqHB6VUOix3DEACDllzZf0Aq3
7rI9MF266t6IhGwbIVLgA0bpr/ejvLF8xP92hDxD9rnbk5tVhmvyZj6gOLsAuJ+3N+xNwclu3GQB
rd6wijas197jRvDwTP9Kdjz21Pa/xAF601o+hf1Z82Q5TexW8bTpjheGPMpIhmLUZ2lLmnIfG1XU
qpxno2FaK+wQNcaHOSntZPOPXyblWZqAK9ZVYgf10463maDyVHZEDW7KAjUbKO7FRa05AIVPFkS0
uMLLDM3ljoslRZjWsBOuTOF24U60VFYj65odvfVKYDedRGp6yOpHreJZUjBKRC8/Z/aZrft9kUx7
7DGdPe2LC9vFKP0mvvNU3uVyxEHRbWOjEz/W8sWQ2dLO+BojLubYIbN47triPLOCUUyvqSbPACDE
LFf7yzW+MOPoOTC35Qleagm2Llz8nAj0lG+P+JI11Sy7VJIaiLp0Sfw3/i+M1QKNqWUUIcg+qcjF
SiRAv+x1bH60M4RIaDLj11OpoLPwvyaPvVLJxHiIRvGruWtZqgX18IM4BUQtrEt149QDXU6MaDn5
NGLvCwRXNP4O8sF8ezDLhRG5Fr/l9qlEu9FywuJGbPI3cUtPqBNzdiMcvHCkCQrpfQBXdZ21uoTl
kdZYDPuBVxE+OjxvhVkgK75dQKgfhcNB5HohA2qKGYYFK6KbSNPdFK62l/XTQpdTqh/ojZGt+Yzf
01NMlojIpBbJhAoLJRriHr30nZiLPGcPONMlWh/6jDH6rhXtWIlKi2ASysTJvv2TjN2lHOXzR58s
rcDSiZByF/N2CaZfOLHlUrp3XKrQUh7y02qZ1cbPGpPGdzgtJx3ZBibet+KaOGHHqelQaNAg9dOo
kY0g3WSnaa9vwvxkPc0B2l44bjKsEb6HisKzAtvN8yWMoyWxHdmoUxAk9RQ04FwGgx/YcnaRUQYv
9Y6i4FFdalGN5BhZyy5RIiMOY4yeQzqhgDupFri6Zf+bchjr+lwmeIYzUxl7qlruPL0d7t1BY+QI
Pz/RX1WKScXzVUlYEWniUlw8RVESuHba//24MtX9o9HImsRyOcTYsFkjSRQnM7+YxOVKaCuOHNpA
myzxADkREfPOqBVZ7bjoGjXKo3Vd0thi3rc3hkyVt8GH4rQNwbZkdC3gqBTahbSHd6GPlNRJqDwZ
N4EMENsH1BFSfp8tLlKOalpPKm/R0mTlmmo3eDpnSW67Odjdj2ETl9UzKUwnmjvueC0ZbdawDPMZ
dAb/xlYmLEkX2JFxgAJUt9A6JmWjWtuMW5LqVFwv8VRmln6+SEHIbX+QZzm6XgYg4rhT158Q+XJU
irlXwlnTscyIJ4s87pXB2QBVyLd683zKZPiV0PDMbGerutDDS9K+AOtDKI6dLZg2Q/gj/MGdpdJT
ceT1hW9foGAfBqkNI22ImL63FYLXsgy/YQxUR+n9h0YkPX3t7C15DrnJMIUKwobP2aDWBdUnm6El
5DvfiAJF6RiIUQq5Nw2LkOyIluY59zE+9D25Ei6gFZVa7ZQTccVbTrkkSr9u4RaXASj2qbr7li4x
KaMna9ksRBVVA5I0rdWVfVPG9/TulznTau3IR9X83jJURTfKze01m6uO8hVMND5utljfL1oVB8Wr
mL70jS7OLlcJICPI5ZiNtMe2ARk+KaSwiEhSbdaRp2BNkwSfatEEqEgkartrj/UcNtN+3qdJ/mqh
SRqapHS8rTosdPKXY0HYTlvxjJBj5FMIZZR+l50IHpvGcHVGCceNNs62TYSsUimVG/PfrtZMj1Al
EWXkrKXU7N2enO06GNQ3U64qfYJOlHQmAdpGaRWcKiC+5ar/RqV+TZCJrvzM4YEvl44Fd7CdyaxI
yMjZ+N6tljJ4wfOxuOw8w2PwWRDf4h9AKG44Ek8OcN8g9vMC0++3Ngdz4kemWkOnDsDMKOjSPul+
/hEn8eB+Xdnksg9/PN2tQ1PPiHDcY/VY5dlBG3rwIHwuKoOOQYFsxZXbjaX/O/1n5429rvik1yDy
NEd9G8pwgMtIjPwH18y2a6FSKE/ChD5YCTAKQmNbrcR6s8I/PX9PVq32tyDV+PP2rNElob9fcR6t
JsZzFhkuxJ8ROQr+GgX857YD9YiraKRGYCwwa71IouGToUdRtfBnkdwPdIOJsajp5v3YPGh6Gegb
HWYbG5+XxopA8m0tGtYvePGj3qEogN8VU7MjiAidS84DxdZhPARA+qnqFzvCc31CvHAEcQAtOm1W
EBlbziEUtUXGn5D98/xkzwFjKeopwRvRs5qRfHJbASaKJENmNfMQ8Y0qNEXqtqEaAT9Q7vaNT0oI
EzYLsbAfNTbHEQ6TIaeleVDvREDcalUmLAItL098yvrFuocMdQnlKPTeBw090rwg5x+hkdBybrdy
LZydZBeNEgQdFBJtsu7umoNSDZLkfLmfgkZc0G7R2Iiu6qMm3M+HCU832Dt2t043SepSEji5xKIw
xFb+bhTm5JP29tl2fHaTSfiKtRkyi3fJq0/TiQ4wsp8n4XO2MxBHvDXrYIvD26c7rVzeuVA5s3Tz
ra6NsDrDLDrAgOgoGsnzWAe++GFqsoAbL5xkH9C1zzCiFsGSn7ofb8jju+tYwfpfq+mMM0KmBXAl
uy459y1nIS4sQ67vKjeh9UNBKeOCe+ejiB/jnpPaJFzwECFGtTMTpzveXNOaQKv5id3DVy8Go9iH
A/O8DisWHi6ko5O3RFaGaykRVj0EiG9BankZ38W0SxWnfAPI4/4hzOH1PiEZtGgA8mnDR5zizY9J
nxbBO9n/NVOkQv8pvFcmFRbXa+2OsQAkKPVb2vxzQEyIGyTI4L6jKF0UYJjzHqVLUvU5Nl5fhPyI
lyaX8L6RYJl8jTmSYJl10ud2ffA81iojSLmPwMiRuzihJnDBnsHNJBgQThW/Sw5uAkVaN2fu1YOP
jRGqbVsMNszepi2AlMbq36vpqcL/hrz9xHgnZQ+JkjFoC6jBciyWtk34rqYGJjkLwNIm57oJCosV
LMNzpXp0lZt94f8pHrXhGGycBmRd/M7uLOJTX1ey7EJ6D3jkB/ohsdlvzu4FRVwbcxJdj5MYVl5M
DGXBvlU3tg7SyYD6zr02lg+bv/ug0gAtFv+DxuBkNsyRLvFUAlDgpDP4GR5P9C48k7L32vMl0ltA
ahneZ233ulUhHuhqFBuA6S/bPQJXBQjshEtdhjk9smoKhwtiTcKLhRt1GW6vEA2uD5bOI4ii00pc
EbrHPLrtZocFgPRCfwr37PB/taNU/BZzDRRIIydQSUo8054hBubp32YlIsXq0xCNrAwV9ri7PpOw
f8XAZ9cG9rwtk9nB5qucy6+HrUC7Tdagb1JJFd8zl4+j9Uec8CD6l+IGiTe3M2iNzzOPTJcmluNn
wDCNzOj6zdIpwQbMVVHsXFw7v2sjRKdR1e7+pKNtujQpAESUlQ2z0AUlnwWyTRymO+efbbWszzkv
b5yK4n4xL5TDR0PiMpdK27jA3ITHWJPxpKbzwDrF9bql4wzYq7g5ksxQtozxe7BJDSCpgNCO8uKB
l8UklnvhqKARD7QGItGUuIgIvId7/4d0TdaDKUW9SSegdqDChOiktwFdP4CTt2IreyYn5vWb4Xel
KLqxzGEe9OgK3CLWj1s34D9+dhkjXvcDiPV7C6NMx+Mltgo726UxcNykUqMuI0wmkLdUJWExXDtm
/tVtMZjEB0NI7VO6ofk4st8NbVHU+7dzWxah1s1v412sgEY4gJti3pr3hUOFDKFXp0SBx4FBkgdc
GYwucqkNWORNEs5kHCrcSTYHVrxNyowLpOH9bpF3Lf9oHJpOFewIFZuai0m5S0d8CKy1Bsr001dv
1dNuAcrogGm3ocHJ9n1V1KUjx3Q+ZdfGoMTS85e3JkViDtgEI5L0mCbGApxMzkYVcH50NCR9ngur
nzYHM4AX/zwhiO+NTNc7QVXqZS72HOv3lSQzANoAJ0t6SM6XzlcdN2b9YJ2kJT4VmoIvHFo9L5Mg
e2payDb2JY1kT2w3PAkpYi+2laJNccakWZW6kmT+i4imzhZjiIQPvCCcnLpKSrXLm0wy3rCEvGVk
MjoD7fG4En0EZ8H56JkRdJxYyHvV37teqfuI5KwlCc5Wj56eIay3UicJHYipxPc0S2PrSC1jwbZ4
9eLVvEKO2Tu5/cB8S5MlThDXuPfwrTGAOhOE11ME5zs+nsW5KD85PDhUBjo5S4HoRB3iRHfoUjQE
S0LShNwOzSPl+LkVQ/0RBf6sVbDAzy9g7fpe3251S7K7G6X5NREnbs2kUe/I4gIUIxeo4Z406UMJ
neOOrfU0rYl9pN94InDVBceFfSGUmrZbU0heChv/35ZQ70EzfAIBDspA43Ovy36Q5ltkTQLmC1Cy
kLDmIg+neuSwIrcfZz8obqH0X2l4oWUxHxExJhfDPNEVLiqbSx0LqoNn/RVQrlqliSXQjKC/QjBV
/gCuzDExh/2fFfMvzKg7VEjanz/k4pR2GJfZwqI7FOFahU5z74EnS/e+3R1cWm6wjL2pEFbi15bj
KF5dc431may+qvG3p/lmvi/lWp0wd99hmlF4vUvlCT39QEKfGxMiI5P5v5Qyqf+COkdKwa7VFMpA
gHvxfsrta11RSEa+PJK9jshME6dgQCDWytgQzKb4LjJJaYDJyG+E9bp1wZSfphqpw43X+XUZ0EYm
X6/YwTBa+a4S6zRghiBspD0FEIOshX/cqHk+HUgfk3yBNjTsmXg0MkTIy1lnyDWXVrH1Na+4OS8K
AAz6urLgEQPJjF5V8AJOEBoB0RNW23x8X1vg4maA8Nb4JPYajC0NHTOLPjhnr6X55MctSZ3keKtQ
cgVpBsPD20UMERahdHHXbaRSBN+Fo57uoCrAF9gtBeq730CzQk2gfvkGSLKaC5VAejpE9iQOL6rw
ymvyeMfpQsDlDHS8bnvkamfWV/G4Ymgaugb/Rp49Wi9SiSy+NgQjZLE/E9UAhMjmF2/1ap1UG+KR
DAC0dtZHaTrS1W1A1D4o7dafkPsNrtLTZnzg/raZ9FURicenyjqY2AFD+OiDQUEKcWkoz/WzdFbn
+J2XDcrf78i6ufz0ZQAIeQbKCQGPNGjniXeDQb38peZZ+Xol5arxM41dyyLehXgRfJAPt1TgVONd
+92zO0CYVk7UrcrwIgf+7XeN2YjBnIUAcJJAWEcy5A6FnIdHm7C/X6YXXC0s2XAvSMwzcZr2Jv2J
ClgJQiDhF2biSb89Rks+LJ24LqwY//kZmhM7ovVTy3yrN6VBwGO5ra+gdzwBbs3dfEJrCtRxeadK
skbMwS1yRb8Xasu3l97Witr6dW2l0tWksJGEEQn1nW4Q/P+xBo0l5O3RTScMfpoZxb10is3jp394
uiOGNVvtXEVxmuPH+1i2L1C/kEywI7LWJEH21iyzADLFVXuaXkyLNAswxkv41RDOXDmjnKLD1iEV
eBDkAAKdNSsAtcSj1Q/Qs1456UDZfJBS/I8RBHDDWTEKIkR1Wj2JiGvC6EDdcyTxJqWiBh3lKOYq
Gu70bfDyNxfnXl1NHVXqsAn9u4XrvUG9jBmIhf9sHcaKg9w4e3fwAFRVnIQSbmJwbeXCaX0rlVtA
LQwmC4K3DFX2WvseT/vEU8r6K2fvuF/NqF0ltxL6wlXsAp2hFlV48cAtWcLMHzXu9G3NHuxVZfAz
LyzgFREeXwho/1VPG+Tnphf1L9SeySs1SBb7rSvDmjQm6ceNTsWSTVO0m3lnZd+rY3AR/cDPiOPM
yVF+MrIM66KpDOG0TcwKFWRbQDSAjoLW68Vh5vokmIgl6Zi232WUt1e0hSQ2sthPcjHAET6Om+go
WihRfYTq2Gpa9RFQbiO6ttSF7L6YPbzRZVeyfDxL7uS3EuIwIZxIywnN3ezPrmvK/wTJXEwG26tu
CApG7becLUepOCFt7nYjZ6aieDOH6OnsE6TRtQRFUpwQz4oqqxlhAXdJnidc2VQIzdS/uYjUl0aV
MkSdYxbcLkdlZ6+Ck7ouPUthEOT6B3h0NjTphp9u2sNzrmd0C6DZSW2kzOkilH/HrBj+j7hfq6ga
6yVrmLcSBg6QIlHAG5RdAle66gTna6FNNjq1skM3vsNaJl/DdSgidZ4RfmXMtxzh/JWSe923xAB+
LN7HRS9JER+ttI5i/RZ/vXfOey+i/GS3LpRkRYls+wMVPg89R/qt28UN8ek+13hGgBSkrqHyXgOz
ScoUfLXkWHZVMD9YLADgRjm46vUMu9PXdbmHZBLi/LhMu1g03rBpauXDkvj2E6pqvFPTxFhValli
qSsILqdWZLt5mo1130esUhQN9pCljd5SE7OUtGpJqWflBVw6DKhKo+o9txjyN1ukwOoP6qldRt/p
i+kzFW0vPYTh30I0Ue+l5S3kR1CE5Q8HHFvEP1yYdnqWlx+WAnZR1EzWRRSi3J8708BXBHgdQdmL
h+iwQPzW5dWjUUU/ShHwXWcbZ8KNhyLLWScBmcM7FdNs2AAeH8F+Fb+Lh5UXQpNWVW+8S4TjLCdJ
+c0HBV9WMXb5FEsY40027aIcf034R83SUVHEr8bceDHxHSGAB6aWEeVcmAziLtqiL+AL7y3+iFVW
VujxJEDCXTHa/ZS6eS+ARQJY7cnC9J3pPvwi3FqQPeVVmzv4xi3GlMUy4wFMaP7Y6aTYzd/EvDfj
kv4dpn7WtHuOcoMufl89896PkAohL2ay3IcY+YgPWZAylEH26TyhKjVHx4T3LP2isaraMh8wMoR3
3YgtIEKUN4pvo5E3x3RVnTD+spwsCR6LPAU6jmCIDsxbp6eBqbRkgk39rtCAnhz0LJ6nu4xWMq4V
7NmmkODcTMeiDZz5xaKFvk5oTVsmMHfQUGPGs8Q9QStkSQ54+oWA9BEP7VeDAdEd6wc2K5m/+OuI
GcHmjuQ8+J64p18iW6OwjBSEGS+3ChdRkb3ivisPKCSNGCGv37a1ZiI8t//eaUbJtIruiuEJ4GfN
fJAFVh/kOP/FUer7QGJUETSLvYyXsHQeDexS+R5pMNsleH/+enTZPwyNyVzK2/zolj7Pb1zKwslT
cV+pMCSAeRUpoezleyic865GZH+Xbwd7Evut+Om9Ej3cFkRBrPs/a7vWgNS0LTdLSDgIiHCNTXHQ
thJgzJEdogdLSMqSJcIcEi0NGpNeA4JWmoR+4rJ7LwM5i8GnFyFJrZXLsz+WGAmFgCcnY4H5nC2h
/lyNt9iVoiP1DdgK9VVUeWBIs0fkfTwFt0/3Y+3bslzav8VlWpar/GeUZBJzWdEETHyD+vbwnXiR
xOPSw6GdiipUf7GP3JwWpnDdiZ+h7yFPzu9xTS3s/Ib0/jh9ohQzvR1EYMbmb92yJN9/xMYWxyAZ
IIjdE4pVwaiauX8ClMnjbZ6DzMl2QCR0aHIZAVFr5N010OnOzV+xmdOTXxDhBjRboF5lRjQVCcvm
aNHkD13s+WYzqOJXgFODMd0phy2BkdRkKV4/3OKuHB85CfYTSIbfRxeEMgC9EUb6IY24lNDiENaN
bci2Bhe3WlTGFBq0J0ATAoqBTUFFSbz3IVpeEcsVL/lef5RO7WFOoY60IkgOycF8v+kRI5wQa3bw
WVZOKvQXWxD6wkLJ/+gHM4A5BPun9eIGt+B27PkpMaEmBNE0WFXXisRUEItHEDsgZ/Fkj7DTBQaq
kCUlnLFr0JoafxbDNpv+EMp4RqaiV2qQqI9N8nATzctjD2p2eWBPGg5u35X3YPHJSGkzciq16Fd4
cp/v6eSYfiBEDevtBHUBPftnmVywBd/tX2uTXlVxQs/wgQ2FWyWl+B+11DsJmVd8wWN+FqtvdiPr
4mkJ3ITbgdrYD89OIuYMkFdV2bq+qAUWzeJRom1x0KpPJ2rjrIkPl2CUUJFQYkEraG164ExOzhxC
Ui3eqMFglL3/C9i0iFEoBDch/tbQg9HkXG+jiYa7Zpsd97SsaRJtQ5xhWsGrxa+irzegHOOf+hcr
EmFHwRdNXkh6Y5UMoUvJkMnVCxU3fd0bEKxk3CHY9qqBAsfvWaoXNkYgYFFWfLW+bcghVTD32dd4
2VSgS5cZRBelwAmcjZaDIFtVf94dhMyCo/3vryKztr0Wokeq/YuJuPuRZHR+4ZdX5MWueAAm3d56
zPiOZikbTdPVHTTyS3+yfviS0FXh5eJVFNrAk+QPyow1xKaL4UqEljOjoBJ99mrNui6H/uUln5cZ
TgJ8JZOkwZKpQh7iDySAXUiTobP/Q/pg4k1V+uYvig+YZQDi5vLmnEYQOFAAQpIdohPj3tV+pGK3
O2lcbstgf9zgGc9wfdEQfMrGOSb6mnCdZdvsd08yEk7ggxQOFHklUihorMlatJy1iVYFe5wnxfuS
1IiFNGlIf9a5uFIFxdb1o0EwZvC0F6zuKxMqDmVCftMeMQ//JZ2T9wikmhWVoHzLazJimSIjWw2B
KIDis5FEj3gkLERlqXN5h3AkaS/A1Hg12GkqAmDcpz4yj/qXjLzuAt3WEzSnwrfLNsmfpN3ENbec
sojPHXMHY3ypZshFrDJoMvXSJ7qO1yK6JRghkBziGjt5vgt7dAi0OTO+I9odsQzO+zTvCRc3rQz7
zmIGYgVjOxxVjxKrnQnoG0c7Tg64LOd/nJUKf02mZgJXf/W+cYUxVG4y1qJ5mEooTozfnTbu5NKI
QP8zh9Vx+ZcTh8OlpvyKFb5iol87Id94zjCOERsZ9wLq1qWsNv6XDG963a3O4dNoNBm2ETeKFib4
6FcQ40yWtXAZlSpPFN51aMQGLiTsUxtFppaqOp059iOtJiUsbRIHFKHxb31YFeV2BOYiY5pGeI64
DUFq75Vpk8gv8rNpCv2eKkzMpyBKDLglYWApqpV8huRiZrlTzaiyl9uiDgF4/ijYTbCKDxaQqiR3
mZxuNPZtKgfRWb0l4HeNRIP/V4QonaJ5jNnukbjdKqSC+jSyGncgWB5eO4jehw19rePAvPsWoLR9
VkIhmTQTVyPVzaOn6VKm7ATLycemby58ut87t6U8g0UXprSlxGqHpZr+7mYfVKT3X0Z8kDXcQWvF
kV8bsQmQ65HX2GbCPW+XskGoDpuZb7lDs7aGInJH7Ze5syb+rl6ARUPw9h8z4J7fiQB9TTnHZTue
6RiyZG41nGBqqrY9BeuswXTUrI99sE2aAb8l27fAlRseHKTiCaqUjACEd375Lv9TBksoSV8EnjL3
An0CCYYHFyOS0beHIS0DB9rLnRRS0GRvLPwriBwOIJGioJ++zT3RRtGPQoP4lAYilVBKbJ/gjyRO
t8oGAkrW4rpf2vJVvIxiBydPn3wFI0ckJr5qF5GVfF5WGrtCYJVBx34mgq4rKA5SsyrfXFluSZvN
geWIqHnTSK3ABj2uJDOnNCY9qcYNPP80FfIHKi2dfLdcR5unirLqUibcoJqq5L1n01Bq5QT5QgnJ
///vkaXZyAS4pTbXIMCwIcyd3x/i3JIq+CtEB+Hi56rLX4RolU2Lt+Vnu3DtzcaPocDJ8XyyaMFu
vSUN6AF3+5RvIV+tiUkY0rrxRwN5RR1QZAijfjLPHpLMtrihMbrsNmocr4EC4qR1V/cp4ks0yB7t
J3Fec0Ip6KgR/hwvLi3HXy70VBAI4jlbHZ4dtvuBdxRM8/8xsarNO5OVPMNYS6samrDH5r/tNWqD
NLDGQXvBieRjkebC+EiWYN8jF1b+W1Sb+N248Xquuvb1U3/EpzR/VXppzSgi4A73Gq2g6HL4ubR3
F/3Y4KZSsw5Llwotzxb4I7NkN29tGwdeHIJi0aJBWZjAq3ynQ6PmEoMZqb5X8kmr4a2iNgdNIlI1
b9qL66dxNbA2ZhwfD8cVg3uogcH8KW4eI8R0DexVeH8hlv+0uh6D2HepoioU+Im2Cw7gQQgP99g3
8j574a2p+YBj7YI//MtAGxQW92XBRit+BBNieDxqRvDU+du8VZng0TykxIhLyenlz8jyfxYq9yfb
q2sgeczilx9blQsh1/79yKYBUIlqjilNbvLDp/fxUyBoFSA1kBmPuizEUOVCf3GFPLEKok1lrumE
NrRDMMbmx8scNcNeQPHGacAl001TnDa4LzzTVjiEwi5KqBbRo6Jv538G/trj0zrNKEkARExr+C+j
rDW7SLKxBfruhBvTs4b1KVoVyNKY0vhzp42gEokGB5XxBkQE+3tvhofQ4e/1UpTSymCXa0Bd25/4
H2Uim8E6Mws6QJfIrPtFTnOE2/PUbyoMetJHbTLh18L0D+lRS7RlsFvbZ0OjKH1vqFDnHPHSBCVl
uyHwpFrlJfzRXmRTm4S3rZW0QxEEe8/OcgMixP2a1xV8KV84dZivxw3c56ns4dHBfU27wNYkRUiw
SW6d2cnEQxBVJKZxIMR/KaVLIOj5auu07JKKIkczK4lGBCNLQdMfp48gqbA5DrVb4rNlwra1HCSr
nxmDmgPzqKOy8tAfALjUgpMHFz3gxiibery1KaaraGiJNMVNSzltgMhnNJggWAu5bE+XfsPmi46m
TYVXkI9taB1eEhCqR0OFnbiVpupJuFxDSwFwSAGAPhrjo1fPPf4EX9VgUjcRHQyFXav4I8ARlhxl
Xexr4tU0mwx5Pjmqie3o+bgPZcQTqcPYv+Z5UmR3e4zsPRZpM7O2OQAFRE5K3ydQamsdCkWbysd/
fqDgBeLTCNTwTCGK2l8mVv0pvyMSxA4f7fXAu/QWOpf3vVtt91GctD6pBad6y90mYnnG8LXCRrtC
3X/8QHkg6KxdA1+5C60Ff6ELGHNJ3eZQn/kr7Bn7q0HFhv/rphSpHiwNwWHsvzrc1th6lluoTbk8
IUIG2JM81oQBkbwdaC1mQj4cKSkaYFxEA5uW/Yk7ZViF18IYo9EZCNl475IxdWeNNaTT7WcdhSRW
uu86Em8EgI/3Ba6ABBAmaefOOCZLfLm3Retq+ErK2zmVa5nucQza8cGN3K9+48OBR5XH4+X3tMWx
Tp5R96NSFb/kA+4hHRYpql6He5HHUBK262uKnnO74ZcL0QpIIeUbTmx01/X/REWYYbecNRvLNgsx
HrXRzriQG8Vd4uOy5qf+8UD0WLN/0A+bdG2i4u16zCuSF9elc/DBHenlWu0DHI0fkGQCRkkFVKaz
yASMcqEBMgCHb6GyR00vKx34BQRjHNWBDXwxBimmqy/dDR6pVblZVpS5DpGEs9YgrxMcb1reKMGq
kSv/dObk0vXprQpiNtPX/vVcmoPeXV/UsbchP01qhH0rOrZcUn8FvH5iqXHDjMyxKR9ouoNg8ZwN
fvdMmusAvgok68RJ8Us1C1/A0ct4XvSfojq4eXYk0XwSXdQLOsnMzFWveXrubP3hHsvZk//7pM2P
yOMcXAu4K67v2PQUrhx4UHramrIGvcNDwKRpBXmtWevjKbgi4pmPDiweTQoWl5b2zGmUMeWV+oFz
6UkIYl5WZWD6SlIcckC6a7T70Xqk2Jklhpag9NmLL1QTtEcq7usnvpyEbVt4V+f+nV8vwl5M32SV
wcM64fll0TusscfqS3KHrKP9DEpRiau46ZfhcRofIH53u61YhJ+q8ZFj+osUOc5ziSRegXE/45/Q
D2a6BL5Hk2J3uNNE+ZEYWVqGfiY6K+2Ylu92iQwr7kY70GUkUOWpn9hv9n9fGSFpOsqsYKudpd5q
wLw/OfNabpJwTQ/hZygPrg8BdDZsVynaXaaLpmMWxjd5rdGHIyIaXMcbBxWR8ZB/jLPDLc2CbLEF
eYL1Vb02UznxTuNxWRA8DNi+6cxvHCPqeaAZY/MWOsERe0O49QdrJP8v1wXxQYlIUj9jrS32GZYp
FKrZHFfW8bA3JctX/fdbuB4KVdosbBhs6R0wASL1qwtgBksOfObX9Rb08WxNnqsbp2jmBcEGeY8B
USozwrq+IN6CanaGdC8nbb/Q0vArB6NGVlTFiLVihy4RVvBUY8ZfI4/6RCQwcGbnPfk3xrjjbleF
qq4t/zKx05bsYUqmsPf8WWAAHe57tcBBbe2Nn9wf/cK8Hf0bzzc+k6sWiqIF7MGjZs5wXvgX56mH
H465j1XzwlOnQkiR9PwtBMBO1XJ7Sp0tPDr+rEz7k3nlsHHyWutAV8suAastlEYyui4sq/SoHxHu
q7e0yDRQK5wXlcrZqAifoX9e6W8JDS/RRKufQy0oAAG43W9AaMpEBACExkj0h+jNhfyyjQNGBCEH
lKmEIXTF6279MsWNb+qO8TWWoQUKpOvXu5WgA2yUHVIpXMImJ3ralJagvcnFvlh8D+FC1OoTmA61
JKBfevaxeT8tPQLA4OQYjOICghEWDi3QK4VB4zsID3BHghXKZO01L4cUwAovPApp4wJlT1O/ZlFH
LIsr9cO4mJRkXsQ1scVQG0ZXOBrkx4cZMACPxV0If1fpxZcwtPuTL9HiuUW+fmqCbV32o0zYfq/m
DTFyF0hQbZerFpByEaOXMMeqFYLCIy0s/gbKIRN6itEmg+3g9BiHkUulxLPElt/ELBi/053SR/eC
B/ghifAAplf77aewfIhr2TORZr2Rrnq8XM15dOzGJKEtf+/QCGBB1cBqtqGuZqicCfSgy0Xr8nwb
OO2YKWObGXkth+p65Xw1PqmYzCLk/eISqj7CYeHts8jXyNkf0cfEu1bbxEkQUbzBHFajCQ1vjWzV
XwBOsL+SYMX2XHsHog/jrzyedrTpV5/WKI1UJYjlZx+JqaoSy4TRaE6fUQkubCYs/ZRqGhbqd+CA
s+mx7tXS6fsO2zEKFOEfF3SazkV0UiIhrlwRmpmFrJWzFFsVMlhVgdSlLchlGUSdWKyx0OIwMskw
Ezsw9YJvRjRncAFnuACwwLc+ndQTgfmr3gIyp0XF0iOGdRYMoUMMQmPzXXhMqTGnjhMA0pj5w3PI
FMAIemyy01lJ//w1JGRICwSD52+UnjELSNReJoKdpkz9I5TuXq8Kl9OHT/7RW7F8voWBKSnyxfPP
T94DidWZ3Gdn/o3pa1xfChckq6ShD46UvX55sWinTpZwUsJNmIpcrk1AQaRTiRQOdAdyJbQcS1a8
LMxz6E+pIBvJfhpB34K26jbpVSgZ+Raw9rfxk2nJqWDPZ75Vcv1IH0XlE1kJMx8oJPCjUliuEUCO
aJqz3/pcHaTPwwl+ok0psy7wFqCc+EwI77MFmGCb5Q5JvPqxaMTzF9g9iUanFzhLTf1TI2G0YwLR
ktM1hSMuEgToKK9UyfC/CKhL1thhTd7yHcvk5havdZufG/krYyuOltEPbZp621HA0qy8g5Qw1u2T
FV80kQ3+sXRLdpcSGfrwBAxM0Kfj3XY6PpVegtwRiOO7QOGR92VVt6w+zcILTm3QyO0ULk6IRLfC
URO2TvuI5FTqYqNw0f4m5gqRS+ZvZq9Kqj6H4nOtwQDWAQ1kPEwvCsjyZDBjaYuQsEluwwWODodC
o9VRyASqQcv6BHc55Opss6sV6nfXN8dF2FY4bCLmnTkhsoG00tSt2q/JHwUPEpgB7I9aNkJW4cLW
xWC2jST3u9I27msE4Q3FlGMUeGvOxOPenhMOmxcVTQRPZjNUzem6aEgAk/ai8Ct8vW5jXm4W+EOc
4oRRqcIYesnMAkCsy9N0sP8qiBd3sAdYQwlc5sPA01cyN/uIFdDgIkdy6UoMw2xJA8qkzwRDysGF
/jJ57R+ICCbyDQHt+i0regKH3gc+qAB6CNUM2b3eJFUVFXCYL5UZvtPwK2cMQvUC3lG78lDMaol5
wyb6sb+VFA5xQ5pyt+fg4mA5pWFRWCFkOqtjO+dcqma9S6Xtt1hVYmWfnmsKser9A2eiL4UgoILk
MCUzTncYAifY9f8/7AqXcxxYmCbslA76vG65Fc4aWzhcFWJMzn4HW8612zRkPUV0Jkp5vNwscor0
2kEsVb2xMlMuNQomnqh91MN5y7wQxqbAsjNK6ZqaTr5xs0fyLTWjn46aQGFVDsWYpzfDdGhrSwIx
NAJa5IQGWHu+eBISib+vzKjZfEhLnVH2CCl/isc/SAdDh3FOSVe+J22Wj2XoEaTid5a3Jd5l9qLp
Gd/8mT5RYkoiHBbOwNNl7l3QLabfrz1JoccPuUmMEo1hDjFXfSS+/50gCvLMZSkV1qwGRRh5fHTI
SqvYaogBh7d/WD61vM8FWo6AnxYali5awXF6e+9jpUNY+/lSX8rIwgNSl9lXTwPyYNCC+SrEYmSN
WFq7/DSbcZGM5BnfI5GwG9YHD11Htuv0jaJhKEl1wWG0w4tOq/PKwdq7XvFSJInniLWt8b0R2DId
zlTO/06ZCcSjba9PGMgHwMg59Ef92n2GvinNxSqSTgfmGO4lxuOUQkpSHqdquzBAsrOu7Oryd1Qo
3F53R4IzTzBQycH7sG5Wf6Y4e6Mx98adAFogb02a6qura8aqYT0L56/nnwK1m/e8CBzOHSmUN4se
XANxrK5zrEW2T34WeIuf4yzZ7wGctwUprhaXwwiSCz9adwjq+ZzdCf3yPjJ3WGSCHkGBGXcHou01
rt+N5nAVQWl6Iof4dH1aFOnd8jz6UuXTKb2CfNn3ppnWcnCbJeKRN2voBI+vMdUMMGn+ibSaZvm+
ylIscRxefSVUXP2Gycj7dStm+mOCOGwCYv0JINhBLipaKGbnZ5nS7eNWjcGsRZHiH0SWZG7Av2/t
u3817ODt4B+7+6wMdt9rUwqIqp22iQPp3cru4wU7Rt2MElLrINwM85BcTtKJ01r8F3j/URr8zk+b
bAjYD0NA3xZoSntZ3U80NCiWGs3TntH21VqeNVCWABLT+sbZMPgS6onV5s8jgLml95jtDzvk2h5u
wiOpA5CCYwipVq/IP9ji3IZVUU6XX2dQ2YnKYLZ31NOLd2+fzc4E1py8B01qmhCCjybH1EHBhWuz
rx4lfrApc6uPVFoDHZnm1Awn0sM9p2mfc8rjCxawLXy3hDe/OZX7L6LoS8cp99SJNZxwsUT0fVMf
6tuio7ZT/qh5Se8tW4NwspN8BSnUBOB/ttHTB+LVhbhxXat9nXD2w/L8zhqLi1QhYgyadxyvE2tD
p58sEz1mssdUJIcJNZyWA7w8QAJabPSuVh23SqnVF4avxEi3lxjePGioBzkOLF74bO8dsRJRbjoY
gGVAXfDrQuUuTj7kdb3daBtRsiAkWlZn+rsrAGUlhsOWa2WfZVgpKeA8s7eJHd0vkPoLnEZEJZol
ZEyg4k7eJh8YbLNTXUx/yqsOLgyyE30Rgw5Sy8vGxg2tdpqBbGSLD67NYDavdC8izcLxotiihlKv
/H2BtDhvkI/1AcE3q6wqJpdY/fZiG1RY4n/pmuMyVRgpCWMuQ9vcoqazBAz/vncRDArSVIvactP7
I77U36eOI/2ODU3eAj7lcHwwPZB53sgVWhO4DdGquBhn9kM38mlriW0LGvgQF0hwc2ASdL2OAPIS
64iu+hy4+hHqH5mf86cUvjSXKf3rSu/Hrz7cZ3nI9/ccnH8sg0LGYr7+qohwUfkYbAmbkIus8pnC
M9WblybG9bUWb8BUW7wVkkTcnSEQk1FWBYqEV6eLuExgNkKgRXNhIuNAnhs8AIbajXGIgKa5VRag
/rSDL3/n64WuP7g5EvOOar/X7MKEDWriQN2KWJEiHAdPVhYubRjEGATbEIRikEI5kj0A/VgRVLU2
ahiKP2vXsP4PLPdqZMhkXUmLO7fBEuqBkz58wmM/LwNgOYcAjF5A3qiW9A48whyb4Q9KcAp/S/7F
EK6gUJS8T7nlPKzdEkuuzr3uaeDob5fKEd0a1Ji45nR4mnlc9AF0Eg+WhwqTUbhMDd48QyYDl3T7
FF5I2ghtDmHYHnd/jbuQpF/d7XbIIkYh1KkYwdO3bCnUAcuMnMKLodJQmgW0QZFWC29A2FR8fgSi
6Rlmwi2e59hXnnzRbLO5WyNTGrU+ucAHOF0Mq8Nlh8BmtOU0mhZ78k91qqO2EwufaYDCFZIxEE0K
BB6AQsLDg37IT25+XBOfAz6w6fiB2BiKxuYHBi67ijokI9s+GHEtm4a68UMU49vheEWGkAaZtP1A
WGcPvs879YcB5zjGlJo2lXCkUgTyvA87l09LyYMwKpyfqgcpFKARf+cgtMnFxDDBdTIZiWp4qt/j
Csa0MDzn9t2Bs1bCZMB39rbW0iAF18SA3eZauejhHFNUD7WAI17sny7PQcb55DQTmWbvNlJxKvox
onQ/Jn8W//L90L8zfShIO69ixtgFDAOkVqQGnZMoDAEsw8TOFnicKM85NrhvGo9Ebfoqk1XxdnhZ
j8UigwD01zrmovmN4PFnU0HNvTC79MOOthcAhsF5m0vo79msaLr4EiA/J6xn6nXQESpKGPZaOWua
Wx9xGybE+eZK1e2CXkd6GGE6y/5TzngS5qnwy48J4cARzYyx1aMrnyvC6Kieox5GhAuA32ggcgfR
EFmu4GI4T4sQ4jaBlz0JL7wUS5sH1qZlA+egh8ORDIkGJt2Im9VrtkzdWYlV0M/FmcKX9myM4hyD
JPwb0s1UnRdiC5Bke8wCIqgenVRVRl4//d5IzOt5nHprewQqWX8YIsA/iJ4gHMJqbG587HWw62Zx
sdvzyOVgAqrlZMJCg8+bXa/hfuGrG4qBZx92Zj1e8Wpf3q59oTGk+fP9d3gtTzED2OUYI4lxYohz
ndswDOZPxdx7mznuvHPn6ZMt3elm3GMTd+MVpLzAZK+MAehmuv0IYjAw6SEpf/JeMMCY1djBx4kp
XmE/DfTLgKp/LTEBhOn9xLeRSt+F42yw6qeqsYfgx1BJPeKy0zmQ90OOIqDTmnz7YlNQ1pybGQot
mI5Vu55pNKSKRlQDe1h2+b2dUtGxO8v7YIFMmq1f9fbQwnOlJcC8/8qF/SFu21KPMpbemBsfhYHZ
i0Nt6SQO5VWzRhxE4BjYV71xMih8EBAYTgjACFiynsRptL2JHNs6b1ayZHMQGrARcpEoZmGarfUy
qqHtC2iiRaXjxafPPP+1g4Cg/ANfymMd6MOMHgxfB8RF2bgEA5AIQTu7ZwG7DyhBeNgnXHPyFy+8
SFfjZ5nc6IOZSF58G8qCRuLpMm1l5VEED+UYfTMEDlD9AlHcF4pgQ3xgszeXLozK5eT/idFYTdW4
AJavxF5Wjmav7NlSUftvjGQ5Rj35ItSb5nFGAXRup3QQKy7fVPfAn6PTtf27DXLP7FlYbCX6y3Dx
NN7B6jAx5qlTYLKE+5ia8BOtMZfYQT0LAhPf4EWP6q/HJ3O4GgYLvNRwUBl+p9dAYSGAr7zpYxVu
GCOoy+MXakDa5/KvlY4OH+7/uHfqlLJcAAnEYeTb3/7gNtMMAcZ8A3xNbrIyEa3uiOCi/3pEfyA/
KTqWkMHdoiTd6t/g20uJ0KY3Fi95Phe2sdjQWi6VKs+4zhRNtnAHOg29ry1PrjVTFBeXIFF+3e9N
f4/DVNUG7QIozljaoC/nhhsen1CIZsh9GTq4kcsDiGNUyh8M2jyxYu27kx65utiT2NCc4YKUdhUT
+cQR9/6cekh2g8uEIksgCqXck5JTeNVouJfXZ6SFcIwIRbliXisd/FiZ+e+N8GbQqG/kf8hRI1lX
P9vGPTKQmTiWLHNoY1hiet//TFr4jermxve7UO33tTQe4hFjrt8/RndSamRymU9fyEqhdmB/76Wy
rnJc8J6o0ueop/FRkzhgL0HPXCUEq5hDuwy5M9F4De3YVVFohPTbi5tFjuiix+mYijGZQQCCR3NR
1g1oobvdmNhgtdK5vpuuLZRunyKTAtNNhL9dHy1/MEOQmS3gow8FYP0OAtnIr71rdnu6J0NkYDlA
xpk4/mfL7yYTmlwcJ8+0Vkjsa2Hs3Io0h5Rj//VX6QX0bX8HqqV/Q5dx3h8OCvp95d5KFEy5XtXP
DZR4DnHk7liuRyTHizcYpUd1e6gVxfAYrR90QAglbrFdI1awXxw84qrF62MnipWSkkQL0Y6d0eay
ecEdBrV0GEK/YXJsECZU1Me9jfY+youS4IjfWtq06myS+b58Xan+nFJTcN5rxvgpkoyIQI3mnQ0C
D/h5xGVgXzMWUzoojPcVjUyiQm8wgX495rEByJvbn9TwutujL5FtMvg6wfE2Wqbxf22+088oyi1U
QF9A2jr6+6aHy7FJc/3TdlMdjrfEHB9hCGuwaskxPjdvYfKzFTzSlcM1sotAPjUT6xJ/j7Np7xkM
4/+y9QtvEyo13wSEABsjnL25QdrGCGYOopHeLpPLW4llZyXp5t5eGXwelwctGXv6tA48/6S+WLFN
Mfl6v8PrbvGj3TGRUshRHKAM8ePoUJOcZBtPIrlYSTPD4gubyybCRv8nKERWiuwGzFpksxV+MKm5
O9kMbvs9GhYP59cOh/BGC3vrt/YSuhHVRrYsl+9q3e0Lfkv0zvLsvWoF+MMFDWoBNqZci1fSnYg0
Dxq6NaFYJgGV08/GcFTmJTtLJoZzhx6dpFTl2hL4hdHdkk7C2V25E5I3GoPuon+LqetKxrI+TPX7
VL63AK2r9AFwA3iKWoAI5TE0q4vY5r/2CrFxt8Qr4AfBA+xFH8wydGZEDsePjTB0eBLT5+71gjUk
NGAc/OJwUUDtYprN5B8dktG3dAjxbqIEsMCzNdrGTHM4Vf6J/I/V1JhiajT7QZJeBBCxDVQTf4Mn
i6bHW+wxunBMs3oSxWsJIS03ahVR4Zxd49+hWcqm3tIh/Kz28uzGHPnG3WIWvNq21fs6YxTREwfa
GnO6a1YyVI1r6ZjaopCMW4D1ZtgYacQIvRsgb3DDfRR+3fI3VTqtZnX2zGEuMuMqBSBqZ+/pxcVv
gaWaxRL57VZwXNlQceIxEWTy7AmKioevbFu/JEJtNioKGjvIk1Ud8MlldG89HIzTlyESJ8V6MsYn
g5U22Of2idUH55rAhNZLMYgvHfndCwiLsjgZSE53QbzUaKXUNx5Wcr2Alv5sBT84nP5MOx2jTQsl
NDm5iNBi2V1G92ubxyGWWrzzutOYY8f8w420zMuOhuRaWiesIn4917q9tCdj9fliB+Uu2qvciPlY
xmvPCJPHLddfxeosyE/GVi8xB5Bu30pWTWgn0fSquqjy1y3xdFqQGGTsNgRGn36kZSrT9a795D2u
TiXTZPuztwoiT8kiBl6sXSGmNFx38q86S/WyRP1ppzb28wz6mpJPHgZ1OQ+84ewn7ncsXp5XD4At
vDn3HS8Nwk5V76I+mjeA3D7EG5XmlcGnup1tgek7m1zzALPgJUf67ehw0VyVh6GcL75IC1k2ne9u
Uujvr8U3lj1EqmlPNF3w/+NK83BwHOaHrzzQcr2FjvC1hLuUYKpQh5slO9WODX/d7ZmHGCcQBSd/
xnk/UmbdMYHDYrvpIWDrDpn0MpZCkbaW9UPHZxgP1hryX9zDv8L5CyJmtwn51X5zEna2z1AGpr+y
QfcUz554V8BnGhVI+WTmoFH4N+HgwvypYHfWjE01VllVXEiVkgkyh8W5KIu0F5rEiclEh+SoYjMV
6De5L+wUZp5ksVk0MA06tM7iUiTFRAKZOalpzx3roAVAtqG9Syv2kpreFhVu0n3IXvgZkrLiEgwa
FEutzysNh9x5BO8/Ak5lDTFbtCAPhq7glduLsLDi6KMeZidWfFajLUwVjIbn5ybeUtmWnZ9/2c51
qOv6+YB5uymeyNX56ncEoCdDSknTbc73WajFEm6HTGeItK5J4WGuSdod7Y6oo8lsVIdivw6Sgm9+
Kyh6tCFQG3JDOEsG4v6gy5iOftooeou4h85l0EUCXW/IIX1mO6pmRaqKHPaPMutS3OT9bO8MkdPc
PQQboNSzQraSyTTxJy0j0nSMj20B7LofYbXQjPOoS2TBJSFxj9cUl/10f9YLKyaocDZktIonAqSJ
1Tnpn8GmNXX5g9qh7s9vJi1o7Y3ahmVitZVGpyylIaoT70w07i78ER5m6zovK376w8XA+nhGOaHQ
Rj9np+idjM9imPpLMnhRjU9FKVUO1PXWY80Im4Yn+NPcRplkDuxu71lOg5MVGTwydn1aNn7+a81j
Y0Fy6op9DBhgZHw6x5v85XSPiywlZjBENJ7U3mTduYJlXeXS5MJOhKH+9S1vkk+Pq+J+vQ6f9Qfh
ftMqmYK5M8FboRYrH+LNw+hKXvnu5lcYeiSoF6jDqqr3JUGaewoiBrCFmAuthkD7OLsseTQZahAo
FbHXhZtoVmf3lGNUkFltpD3uG2LYWnhAVa1gVZcYXYILSP0HtjIm52EB0swH5wrdn7AMo1TlWaqm
GZPB9nXe3YeNY95XChxzFJGlOOW+c8hHRVnL668tRC4WMp+d2t5OS8bPBHAFKKRLBrld5B6EatTA
CEXwVRLSylkZb+h3a27yphahxiKyx/s8A7YoPbsDZnLdgpvx8y1wbwnBIJGZtw6XKympacq3oGDn
ZDluS7csaLShwhQ2Y3i3oQBGteXlT4nGu2tXyovmWQ8WfxcoX3bw+2xtS+P/nU1FwgPOmf6vh/wj
AX3pbXiRRQlwAbciOd2zEfDdXBxA6mgmdlvq4dlqfyhvL72mH4ERCaUC6s/G8GWYZK0BhrKj12Hi
36RUcVi8k/an1FValyqqDs3RixFgwlsqTskbLNdJr/USfZusP/X3y8JnV+TAEqWe1Yr1AcMLkU+O
eC8ast7qJOirQRcFQLfNMiWbhPp/4wb816PXIiFgNtG9kBjKs8iIAitaY4vhEmHMGhLFPMXQ65uM
o3H/MYxKcqwdCIF2maBNuIDIWVwnstfk64mwV4WMrE0jNvRHi64lXOV6nESWqTo+AFt0C6Pgdxll
CAzOj2fBd38AMY3sHZrJ8TOVYcU459Kfi1U2wZSi8Xpg5JsTPfHdXUtqf94URz823Qlc3J7LnUd5
48M9XnA2la1eJkiUWjG9BGk84pYbS9WNWxTQcwylzkoIWVfRKZwa55I9SWgP8r/Qzo8N83fJM10o
1IlkOa9nO8/TU5Z37aLKs7/xvZHkT1db4zWrHylBgkvJo2SOLViHfB6AATWXV0ClyXW+qwpzNlYJ
k9su44LJIQzDwxCQ0Nn4TCWKa/TkXr3FpxmpO7RREw79uDuQpkyXTkFX6IYxG3jgo4Y9silmfTIA
/fYUGgwcprD+KQj35+JshRgxE2Syw2/hTHKkCJYueS88F+EJ558qbIzDsPmxUCWwEsa3XYPdpCUp
zvixA5PO0H37cGNyeyP3DSH+c1zVUEfUMgd0mbYF1E0gclBNCdCWQMQ1nqLi7i5DgWEV0z6u1YL2
ZgHNklPGDpMqbsMBKZkQvLl/28xehWU8Ojb0mpcoxqwfedUdA2qauBariABxgmhq/NCKhKN0hhdv
B7Dgyx2/67SuK9E4ecJnnuZGXmEwf9GAbAQIvBP4uEWb4gWUo4WYpLWQiHplAFCJMMTouQFOKK+V
OHq3zew8zKlG0Wiy1+4TV2Us6GKOD+sUcrVSujxPSclNg7uA0kIod6NfuM1Fwxicor89Dt59o9i8
hWJwc2gyD9vJnA5MgPZrJ2YHpGaR10yB29xGnuveoqfcZlUu8T4Ypo8szm3phwbPlJ1dIKiVc9dY
LgtVkx2fO3cvgl3CEeFWXymO12oupHZ7AlPgAnstv0lucj8TT5hc/XaW4vRcEJO14eh9kZAvbaZU
ZeVcObJ3/O2YXZjgBYp0IENJYZnQ0EEJ3DM1k4FPXlgJoUWAHIi0SLbJAkB+J04ii++7AH51Lh9v
MEssDFWxEQs6Ln9hwYq9YKlQehVm8M9UJOQD9UQhGH/cBMDlc6oEDRWGHVdTOKeBZCMhiKqvpGdk
D3kFUQiyqQEuuUEdSGZPn5OzjIdwGHSxUcgMA9uGKEJd1QhZv9LWMlfRuwdY9N/kdbPbSp6QoIAO
v81WskxovqDUIpyGwKS/N6x9CCcj0ry3wacwMxOBZ/GL3K0a6o8R9xKuchkvuc2p8gdNKyD2DRs4
WoApsaSPeXDTfa0edouM2sqs8w26b3KZ4SHRunYBeIR+Ww3o02FUEN1+icpkhXV0C+zFi/bQDmUF
FNq1uXlXpEFrVUMTtvl2vr44qsaLIIHM9OtHik9nytr5b+TgLTh3P11mcEgorvot4Uhzotr68uAf
0dFTm1btuf1sEe/bZYG2vnRR3fwnfuvt4m07jxJ1WZfEap2NikFZ3l6zqqbsivXLVSONsYTzHQ5W
flG1CLhue7+btRIDB5EYClJosjT9VhSzHZNy31H9n+c3wvqheaIhtRYh/35+r/UsB3OowW+Geyr4
lPetjTtrPhLseyclk/do87MAsXvbDbvW79vP0o5270j97XYyI/PML2puvwM+p7AG3Hy/AWhvz6al
cRLydjoIMQf+ehszT/eq31h7bQ3fLybppx6jFWcDOVHgZaJg5vMow76vDHXjn7Wf0Cn6x0I0fxME
tEO3pSTGC1j0EqQJ3DXMlQ9YIWM3SnM5eJTmOjdcvYphe/KOGNuGwMEG11QrQNN0UK9ap3XluCLH
A5oZ7G6/e6VjFvx5stexTAyUg4zE2tFppZ+SHrlAL0QvKKw8HRoSStdtvMA6vKhS1wKa06l9B1aG
+7rXoCJZEEyw7VHofRh17gIJCoE93HzACvyesITSbXuSGdVUT42yhS8cekdqMrup7Ny+fwRGMCgu
apgcICS6XzVLtLmMrvoTA6MAkgSkusQbl5C4ceFi4lCd9CnsbrpdqfWLFWFO9U0IhJgg6PF5VKSU
vsPNQ7mG6hf5sJ458W+AudHm/H0J4lOuHEMM5pVgtZ47UfUHz3uxlC8fm7MKAxtprsALSz3CHcc2
2wJ2tzDhUIdh98MRC/7D236q2pMFC9maarGCy4n8x6j33/TCdQI0r4uP9eg2z3Eb8LrCKT+/h3lN
7KdFT9ETXTo1veBBKsJU49o4VWlS0BPSwmBzuUTV/p5wCEwVKvnoCngiIc7jjauZ1+mUzT96cmM3
O58/Gm/mYnwlLlTnk1CihauwW0UevoXtUlyT02zFrC/duiyYNbUs0bB6TwlmRE3AfdPD4Xiz4llD
tAMFrcFYnck57HW+uS7e86R3y7ho3zOVP4zJ7s3++wSxxzBDDZAMevN+pLt+UYfDuc1rq0vpvO5Y
Yo0aTNez5S985st5dU5+ohCT25fgFVdUbaPzsTt21zFYfIbkTF5lnS754LkM4skJsdRa71ZPrqgW
t8JZErWdSAyzT1lawtS3WgdcqRRR/gQCAqMQh2GZhpZ33iRJuQPsIqijWeA0Cn7py964FEPAZHG8
tIvPtv89lLj/COy4rudif7ITJG35MtRezIdC3BdYkE5HGXw5JhXt9+G2JqmUXhY9/gVRFNvEE1m/
8nc/i1JKQm/bbasS8BrnvFgiD9T5Vm0w/4y/lcESy6TAlaxA+BNZGOPDAMCY9gABgb1Zana36io7
1s0QGx84gEBTOodGQmTs2nFh4XNRuuHVje4v1oK1kwroS3hEPvay40lCeFUFW4FWEqhZuQHwAS28
RLUL8Ahof+Uyp6vEmbmL5o53PWfABzLwwth5pOfvnDqLcAxGl4rGKw3Nlsi062zRG3b1/akT90D/
dS9vYSmeZgr6CFIVab6Fx8ppgPAu42mslOHuzSWFyIYhgO2g7ItGeCp4686bhvtkJwTDgJ8GGfXa
R6ejxUgOxkLVM9VxkE+TGc2uw86dKLVXCF0ZyEMeEpYN4Q/Us3r7EfbrgJ/txGZ2U+UjRCKRlTrt
/wRiK1z+KoPH6o0eBhuN3g8Of9xg30XvfadA6zTHWiOxkUeFa2NozhpMwhvQVjK/m+aFvuF7WZcM
qvTwatFla02drs8KPG9G952eWCVTKrdHdl2rvQhCAxqhtzUrrgdcdJiM9CVjjh6RWbLI+jxYL+cZ
pS5qk2yGXHptexa8paiyzB1moJtsVqJLigqBXCq+t9lUnLQdnsAF+6LCE3RcBVRh1chZxaJFvn0B
57Bh5ealzEnVMPOMzrc/zqcq5yUohpde3CgWElx8w9rGOgrbRTLFqdgiP7eULc0Ag4/gXwuzxvsa
e/IkpqkB/sgxA/2Xr/45V30bAkzwpGdQbkF4XZUHh57JkjBw4jPI0mvU2jWhKO3vOudyn2PD/P4F
C4fN0LXhCbDAB+81v7MfjvEx5pFbyGpqBWpr9tRC+axJ9VGYVBdHieEnK6fy8SSNVqLvt9qh411H
lCsg4S9UdDHItsQj9HxefqcJDqmXxzhaCBDKiMezldbcwklz2AKB16e8s2+Xt5qLAaPJ43c2YH8s
Ud+krj8A2euvvXRkF778ibh89i7xsmSSUbGmpGaNi2U3bMsGfRHFPEl53gjRpF858SJ7l7wWW2mE
yOMMMSmkuLiooiLs8X7/c5hVgFvIBgg91dNyF7iSSQVBB0pB72fp9y1FncBusUac+IOFX4aaUN2E
IP9IxIHs9okvaxe2PfnU4GFdDS25CRi98/ovspCdz2fsDsY4tUs/+1sup5mraglvh/erXN5ORukR
dqSvUgjXoTstG5bttc8yrFvdjgzPsXjCHFODfyudmgNAWniRtlIBdnEBr85taQo1olHmHQWF/7b4
QDlGMK62O4+8TiYDNwzpbHOcaBrF+3mmXOkMcxzhSf1oVZxsrcd/nCGwOVd4blludneQ8WVif2/V
DTzVWghQLRYviHfSesGoSDCBydNqwCiVEFa6+H6uEDINDvJycO+516ZCvu0NbZr56N0/l8dHFdGg
G0tnjnzSxZTb/D/ZHE+HgJS16nUk6zqyVAAGib0EYbheEziUVOWRbGG3mjjwIe4sold2ai2ThSmB
vvQDyWQL2F6jKPeGiUgTSIUhF1J6HBK+KNKnSd3pLrRbc3j89AVoVO1E2xggQWWHhuoX2KToY8jk
d3mKdr0PE2p+L1k6v0npBbdtvB6eoyhNS2eMpIvmfdce7AB0PTrk9KcYDaje0paXdURS7ugB9zMK
/wNCsoD0/BaretQm0UV7+q/HRMYNFphoSJAlip3FmWtObjRmj8rBrhlnY309OamPE52L5nJmPdZM
twyeJ6bWhkDhGSUCE07VmL9Hesw1kz81e3KbTF9j12faefczKJTquupCthSKxqchgECXoVYWbiRU
L3ilj6Y0ZpJGpiWry5ooUonyWgTlziW2lYiabuM8pTL9YLXtByCajYlKWyTwHIGEhW3DWS6hxfQp
+E8PvA1AbBxU7RqJSqIUpTAqnQyHesYM0Q5uIhdhmBGsqBHYAf2SDKJFXOjc0DOhTH8rGDwNsoK/
+v/GIDhadd+XzY6FywvnLkeNS7+mlNK8A8IHD5J/Cn6+5udj7Tcv/aeWv7hua01ryZQUva8S9L6Q
6xyPKEV259xtxiaUprO/QsnZVM3pi0os9YDVmT5QzAgSMG2iokFqJArWrh0QAEjRAoBhW58nnqHB
AWgAGjECEWrzttK8HOdVL8HlP57x2zNXR1QQqOXN+elDdMwApLWDzNYYrfd013BwoELZk8JkyMnl
WhyFXBsUkYwWzliFNhKJqVvCdq+9s8v3JrSkKBCHClT4VPQKGGEXCWPt275mmItZcxYLPaxA4Rxg
bb6+cK/oC2BoG+dwGI2v5S7Sg+viB2HDwFpVKKTbeS2t9OQGv5I+XpMR0Rgd+1jBVLJ89DBfgXeX
Sn9A5bl05G1ZZSXBnKKLzC9PTyZ1qsGoW8ou1fIQ1HKWp5qUEr+XmkgnPPJmfftmyQYgvWEHKWOX
vQTwyE9IWvyhMOQF+xP1LsMVobHSnbIYOqS9mlotYIaDGYfgufgsSJijSFNYB/Epj2lzoZq926YW
3kfdwdUMTXqvYchlg60CSZYb0jTMsw2j406sOFPoy58XyBtSrxDJudSErRHLtXIYfF//OaiWUCTB
H1br06Dgr7IYohs1ahdzVwD1Z7LQdTk/FbOwZGDiz/Cwl69QPhZMLd/EnEVKz7nJpQT1l3cexJwg
PFCd2+MqxB2psWtVP1LCUCNz1jO3CGLVqwU1UmMR8cLQPWKavPQwUaPPnFNKQyUPwNsPypki4Z7h
WO+uLb0bZG5RK/TAfIe8FDfk3Q5nAVCKnI+Mgbg17uSY5mZnRLnblGIJVGs2wrl3iXUv5pGHN+6h
/fi3cHDAmrYAEIcHs8TrbfnXtS9O43LUlFh5oOXag3iSX3FAdlO5EfsDU6IidL6gT1yaSeK6hnzo
F8VshGWpE2kZ2TkqTrPSbWmhbgISancfYIx2cbSdppSeEsydoDnnreRIutwmHuIKDO2Y1gerAWAu
S/+2rzC3wcAXHELJKZXJhx3KNzCGW4ef8XNpVcneDt1/+WlidJRK3/XzZ4pOBFJ4ld/ItfMAco3K
0x8N+ZnP+JVgYB2JcyPEjkWSi7seMz3BCB7YEvm337WUrXfR1NLOWFL07LD6nMSLHqzAObADXxCR
Bd/IbOISKmluwYH4G9TJXpYXDVNNzAPly/rAPVbR+iMsjZoqFx83gcEOfF8xQ6GtTqc8kO2+weQI
91tNUBdb5fJLi+8uoBXeKWTsOuB9MFvjKeRrYAG4bK+h+i7z17viqVSbVzY2n3kxJbM8cEbJqKl+
qaBZCsV9+ED5XEzmS3Z6CaezHnPxFBQ0qlbeMBWFERVnXwYwdj8Vz2pz9KpDzstcr5rR5Zdfi4xz
WeSmkipEIPoyBaTa+eoTYIo7mTNoqbNH+PL1bXHA+Cadp2pK/ObhEklKtUOSZdOWzFIpy5NE0h5b
eFV+f323yHtLXSpFenoMlps89ll7/euiOKjQD3BNYeguwbZkGMOkI4AV4QJyG9q9zG/asEWRsSUJ
KHlv70gwqLbO7iUpQ2x6OVqPRwqh9C+Ga6A9UrYy4jWVZWTWT/GFqI4nFxX4J3I2BiPdxuKOad8I
PyBLr+IuIQCx4F4uNBh0h+3ogPjv8z8wY6sri8XTBSwnoC3bLJspkrY68RiM40ogCM8pBJIojnZT
tireEQBl8n0xPSsUyWNP+2xiu9jPIq3MexQ58tl07dpArhc5h9bCJEFYCz8N7tVScllgC8A72qnM
la3TDRhn1WHEFkH/qb9AixMnFIbzcWL8k93pjc3F+8tFu78NJDt3BnoC9Vlu0avUfxKEYDEB4Ian
1BJoHDNYE0giSsjADUpmIq6UnS185gHIsd/HuTGGwISoh2q5zp5NEYewEhjyA4u4Ylo7tBMNFg26
lRS9lTliPKcGAEnZYsJA3LlYYU6PsPR+Vcv/WdQZkAdhlGKs9BEg3oDf+U9loxTSj2/58p//Yw75
IaxAD+d86NKTfi4NDVpABEVa6Dikymq/ZQpnl2K81XE5HPYgz7owvHG3RiwYUy2/GDlH1cfDaj+A
ga89vpGoIgGnr6KERqCLAQKezqND77PR7fOF7iVqmuDL1FndwpfUCN/IuHnYLZzER2rQkc/XuDU/
W+mjoELRPOmqCkLG6ZFWkoZnRZuOGkygcgKx+tNIVn3obVGkVLRzEuCrVsdB/Zu5PrrdDGvjoeh5
HkYVx5PLG8TZXFz0kSkf7Wk0kWxtIv2htBIfDKaQTFO0RFpImF/YSHMU82NI3658ZO4Bz5xaHK4Y
LqaXzrDAB6bh3UcMzjiZi0k2v0o/C8I7eB4M7yvZ2fh+hQRDBWLI0iysUnj45vTeupBt4+ab5z2o
TYJr5/RUYJsEFgrNTPbT1uocXKlJE1v0/Dtia6ou3+cufVzg4BglluvSMM+C0mS//Tt2uqK3dUWx
RgtqdJTIQ1iZKaGtzxwjgaDy80Kis+v17I0Mad/S+Zas0iELAVwpSxGNT1DUIzmVrVUQ5m2vTD48
FenvgKlE9WGV+L0ph7YTN/CaiBAgqBnUzTLGbGIzzmv/5qDLiCOnSyrzxlih9fNGv/eUNREDLJuN
SStxB5n2JRqg8LIeVsCnz/gsm5ez4R93JxB5vAGzk39Ek7nA2KMjuHTS+lo0yAC++lncpUTNtv8U
Yla1DZ5JJhuJ/mAh2zZTJ9+XQz2PR1LMDiyN6gvoCPsVvMyg8RMYTaimQy385daR5nqwzP+aG89u
TkOx0RZKrCMkQJVH6VPVW6Z4DURIb36n1EN2+LasQXn4dZdQ9qH7DVHtLRPILBkaw+UbTZXuabjq
B6oXwPppkxtnmStGuVmm40i3Pj1bmciVluWLrJgktLG+POfpRQ8Jn7lu3olcDja484lChKtQZz89
RaY2HzsnWQ24XPmBraJ5vN6ZALuf+ehriS4ZIJ+r063NBSjpT20vFxFWzwAw7vjPAC9hl9WCmNpo
bWsTO7ixYGhLPkcWDa5LnNPhPrhB0sVbWMi5HtF6A4G/uKF9DNl0xKi9GZbLOK7vkznBsP6753X5
NZ0+k8RSmkZ0nNJ700m4kEUhS4UjJWeEPswl0w3s8bC0gPcNtpB8nZ83ElEUbufRkjGsmLESQH3J
1Yk7lFlnmYyInsILnWqE1yPUfT9n5taBVLw9MtFor92Eq+sHKTxTPPjBb6QOXg69ZRr39PoOoEAm
B6uDYTB7y7+q+Q4ZGMKvC5Vu+bcm9GgIUunt2t7Jv2CKaaqFaEGGdCoBt9achWqIVTatUuKT88Lo
3GZG8qADFR411gKxqfvqUCmpTztjzsl3mAutgL8zB7xGCvjqQmsQwuhudKWzv0Y/KHseJ0D3sWtA
t5hQ8403wYFMH4BIXIFKkZkk3fXODfX4quyDi5rLopcAXENoEMmHQPJr9vTH4eHehrMNV7fM1jkt
JLEOc4+IB8+ozMJp+e0na822MOcVVCoonMk+9w+/KgPgb5j9oh4lcTTmC63eg2OEGzXkBfZHgjo6
l1YQC0eHMNJuSj7W/9DX2+oBvtQUeMT0nI7Y2O3ZivEsCZjODG2fIIu9ml9Og4vjyoJECWO4z2Tf
nGfa8nzZiJSOtedY7+O4k4jYmKRKnoVDiMylND9D2GHnpi7rirER3dz342oAP8vwOFlgn/+gxx3j
vDAeDySATmyX4zzbvBykB5+JsxGnlOjeOF7HiJloCtgXsDaODy4vffUnF4yTtZ1Z6RyVbtRhFnsj
XEvbbRQwyh1VTMLFeWSM2IBuRNu8ERS9acYufcVDio6/QUlE+GyVSvUCgzhueDEEna8XN9myDhQS
T9n5nZ7H/tIDmHqRy9YFhHRdVJwI7cdwmLlT0tKCE4dKzpIGs7NdYrgsgQ0YB+K1Ogb5Fyx5pQcu
ULYxNr88CJ1uMMA9FMaKWoolQO+/UXoENUAC2vZrYItIBMMgGNoY1lx005WgbDsDamUPFpB6hOZE
2ZP6/ysgHFie3CBkQjJjT6MPDLl5bNsFy2C+/nR+D7WW2kR2xkyX0FiuMuENCJGukGOLYOwHXuWl
58cLWSZdVrZ+h8WjEtQLUzkO6PlpWvZK1WVwsjnUJRJq3EU2Bsc4MXW5y0quYM4uyCnYNbKAnMco
Q05Akhk5m9ujrP3Z1zY9JNAmyX2YeeBKOtUHLzQOmNb3Jt2idq+1rTqswpwPikmQvH04T1RCNKip
LQR14m2tK7eNvS6UZV6jsX0YuTWizxFj7jnJFRcdjc47cI9NQc4XXKILosVHvqqkClCNcthtnc70
D9SajtG3tgTYRzV9zP9wJ3VLZZobgjJXkN2VC4WswLIW8SRIZ38B28ZVLWita6w8CtU56Z0yu830
oq1/cn8hDzC4azQ52008cbVy7aUIoYf0j2+h3Q7wyIq0Hwkw+I1QqcWtF0jzTirNwiOA4pKN6zzL
cWSyge5MTnzdHgtvTCSe3kxewjCazWzbDWH2CpcGvMaSEyGSbcCd2cw1ltKdRwVENKfoig7vHhvv
O9A+8Q+Jf6XW5Y1osTS8hkrNMB6kJLhjpsMP5IzOc9VNDfXzztwJ/fbQluz8mjFKFNVpIUZ6fhGf
dVSb7z56wR7AaIp/e5qMS9LPrUKt61pDH0iPw6s+oQf6+3zo7ivp2Uxn+oHEGQ9vbszMcTCaklK/
4Hffpic0xMysu34GFe2tWvaIoDxbvnhm4VJtTQS9huK9xwLkR4ZFcE/6m/TWrMtNjqbbKfIkOdD+
rLoXLHqbZu66/NB8qdYcz3+BU+XzD91qjUg8ZVmIOZTxL5Lsc2N+drKhiI18VGv8t6UXSF1UhgFL
iO4L6q9urlOVEFLHEXeao3+7xBL2DvU8JNWaEBqd7/tTzBfQi/rLqbAxi3ggioVdayqvVrqpcw7O
RndNEI2iYX4KeIYHw33GXxg9ZghClQVPr/O4Uvxt4Y0NwSc31KKC40SQiwFOskWuEBauQvhNibGC
nXmoZFqdsrRVK+or1KLZdgTykGS10oIH/Bl9xK/OS37uRR40NaMAfX5382qh8w6iM4KnGn52UoxM
M9cIJMSZQAO+FSsx43ENgmEq0tawkZDinvfA5Gdi58GZz9egXqNKflzu2aIRaVZ/72xXwxNmbmYP
8VeHb7A4r7EM5oUCGUwg7lcTsKdhok++BqimXtBuI2KcFuBFrornsRXMvnosh7Gp7C685QmYObkm
VyoLa4SrMXNoRG9T71RfSzxlE9vTr8ArwB7Xt/FalJaDV8r3pTmiGuTy+FfGXoBx9hw8hybwSinC
TE07MChCP4eqAFiRCUOHtLgdX2WnbNccYDsL9Gi3ECmpd/swLIvUqobaTgZNQtBAacC5iHJzXnRS
hdjBtGMVCpk7CLO0XqNm9t0TlbjjlKHgCBgpHOOv21tzNntIo9rYWt2xunFjYkEawwHM2OOIv7/n
28pLzW+d58m/pt45YMXzNlbstoLmmrjcNDfJYemXPGXT3wd5ml6st7R6V9jNb8SEudunOfBNqe/y
ou8hEYAfgwFL7koJr5lIVWxbQttAM+YJAnuW86Knvgh3MXQsR3ygDAXwLTiX+A3mqAVdkhdYCDWY
MreYGyGmvlXDdZ5pOGMeCXweWSZ4f0f5tDCMBhWvOUkR8LUHNmlhBwGWlpsPY3BM0OeHxB4VTKnx
q5lUX+dUeI0Kd2QiYtRoH0G+WnAnL3hBPC3E39TOHVjssn+TUsge1BiaG6TE/yTuK07SjndlheH5
l6LoKcEBx/xso41V6gwaCT1dfQRxTJUpOglYksJ6t8Phs8n9uzvSTzlpa6fIIxAqmKV/IusCfoES
Pp5TWmcZ0kn6ILr7laU1FNqFbFSxH6cQDgTejlGLZqhvROaLkPlP/Xb0uqjMq/PS7JOlyj046lFP
bTa8eBWtasHKSjNh18K0ME1q85cll4EVKRFpEhieGWQK2zLTHFy4BmLaMFZZa35eXy/M+J4dw2mm
7QdGl3uxN9QvHsEeB+wohdrf2PISQYT6g+eiW6V9mlppNzoy+5pO+r2xmGYzFA1AVnnPOTB6AaIo
yvphg70+Hp7UeQEY9o+FkUFVMoycQyGp52t/p9MmN1NkQ8M1EOz3/w2UDTQyr4karUivoMFv3e6q
TetzRaxhOcFWtwOThFAE9xBpC8AgB4XSlJ+tO+AtRIR6xZbRUX2ha+MRcjfT8WVMT83fmssQBBJw
n0mf+5xo+REU42fSlSEf2bo6JG3O64DcK8/CXcbj4o9xJoQ6XquO83JLkHiJwSC7E384MnDoGvKZ
D6wiWZYcvJFvA9XpmTYGkS61Prq2GVvHyybqjTPOXO89I/PkIKyu1Ti/0B5tRFyfQFWMShYqjBeA
k1PTN7XS2GRPjJLakGQL2uuWxXRQJzun/xuWkHQ/J7fkB4eiiJtlIN5H/9RXjtcZGFT83x8I5kGX
bn+1KQfqduj88gV0GNTK5MD/UXCMRKNUghsAOErjXbt6CCFAPdk4oQKLe16di6S4jNFg7HQxhfjH
yBSqWCK/RA5QIgNAlD4NuY8+rTSfzekT6GRkkdIiWkN8olcvd8ka3aE/efBfoF9O3U+BndrCwrlr
xdkUkRrL013gnn0jzM6cs7FKD810RvATbVIYCncx3GOeOsk3+f65iiCb3lwyNxU0sp3+XZgE5dc+
5YqVpqXb4Oc1z8vbgTC49581YXaI4rLBoT8UXyLnObIqk4zWiyU8MxjIUS1yPVX96G1zYaIMgp18
XYSD3QCEt3lZZvvZslHvtqVFuGi/QXFs64xdNhw8C42hvKmJMxrO0s1iyHMLWOQt1Z+kzpmKpcmh
l2OK0VE/AKhbONSel9ViJJlkQ4NLrMqnYYVf0OvMdfSCdBQE7XK+v53R5C4cznSXnWSWMu59sx9r
iKf4VoYYIS2v36vySLpAmB0CtTig/GDeJfM6ufSZlV0uOqcyv+k2VAFW7N0TQn3F/qTzvDi94dpT
XewsLMoTbbLqE+289tP3Vub3TQbaqKfTpRGidHQ2IIkyoIUZ6CMRFzzuNmKhF3y1Ijgt4A3RHPgM
3GJgRGB2bMrBIIbhaLm09ubuN8I67Cqzg+TAukW7V+0PHrTsd3yKuq4NgANZ3p04towKojvWaDK4
3EeV/rdLshmg5UF1wjj8cAVBNRy+ERYixOTQdi9+tezu2fI39lEvJO0XVeq3IeeJah+kXUTzmO2t
kdtPW9XZX5eTOIVesrlX8p8gi2Zqfap4J2cPuXqdWi8yOU4vT4xsHGjzHcWwbOA3nHjkvcojbmnc
byYKw7GujB0/6fiY7OfIh3hsEXvlzJQVaZ7FYJXc0x7rnek25EpxEMKvHFb8AhnIx1H5k5uyw4uU
3LrjDNpED2ZEE+hy74fom+43E+6h3HO8YB+QgtuWCVJX1oaw2eM5K1jUmYINM7IA2XsUOcEHAeEt
zn3DPpRzMNMTxKvuN3wZSkmYeSM8CfgfECy4CgLAacTkP++FXkaRETBORaRTwmp8BVrlcr2C39RB
8C7Qe9t+Wn4GsoBY76dtLTmdtKXRtpig4B+mWc1qlgKW1+iM/UFSTVieNax066nhWnqj/Sb+sP4I
eSJdMKJfEAlLOB9V4PBcIC+JJfxP0Sho0r4PT5NrWNmxe33yGglMstXboAiABCscrKQDmOA0yyy+
NLdKk5PAmdHyhMkdEyi5tx0Vd9A6cq/LaKqoztQPqv4bCY/oLA6Pk8xGuiTOtRI9Wo/r/12jFkPn
QYctCjzrKpfQdMIlunu9aXb0HZQtMEWtekxsKe4l9p22s6Ee5BcTkBbNHZ9R662oXVGG+vpSh1HI
D3f7Y5n4JkiOm3f61T6jOUhsVVZs2Ps89WzWrXxHmYZJyauU85HgoypICuO2gCQptZwUdaWOEzYw
+w8p8Sf37LYJgtaGRQCKTBNCAGeCfDnBDt8KQ0I8HPdjRVIt0BrvCjTJcYSdsfkFsZhEGTmGwlVM
jHYWu8pmWpggrnjiGND4Ls07mJ4qMmMMnCl/ltb2W6RkNZE44DczznnetpRhFAJ+OYxM9hVXlyyf
+C3hbHzqNlX6Qf8SgyHl7HuVJBHroGinHQLrJex7dW6FVPBzhc6lUwAra4fFsv3sMe6QBy3P8pFW
J/FqRViWhgLpnZXo/rowunJJCJgvDT4vupETJR+msY3DKjVqGb9jbfxMIAMDdwJMhi3CF27bUrei
NG8kZVVC+Lk4BihWl6s2gI7FdE7FconlG7uuue7rGWIkQo0yPO82CxbpG1EFuMdBczr0EtSCIPZa
2jkYSmUyNYDcNtxFrY8fltkpLdQMrU4Wye9g5MPeFMgAfOe+xZid0PyAaTMudQDfTSsXo23HfpQg
xh/mamqUfuC6cIijWH69l/MwgnYjqc3vuR6v+UekjjKfkH3gm+rdSEtq5SZshnmXhGgEXwTCu2AK
ZXfLSyr5LXVpCpRX/El4yUgbEjg8ZJcvhaFQPVShJK/vme8oaX6s0we97WMQ1V6JYMNwh6CAsojX
rwPdhPLOXZs6+6j8PjmKx39tzyiJog8U2dB1piKR1X7h8tdIz/o9BjnAAUDpZkWcadBSYP+1q1BA
Hww9LDHbGpbLOPfTnYXvbpXoj2/1A66y778qV1d6/NA1yyAvqdKVE242yVQ33nJitJa9STUITqo6
wADPeG21/O/T1o9DMD3rG54E+BfmYy64GqutRFxfV6dUuXBqbLjDMSDPp/jAG9G4UmsbMkn6KKGl
Y+hyFX7Tdfzwf4dBrHS9r/HQ8AAkfAt37WZZWKTL6eqd89Ai1KwKfaKF2sk4ws1VGzTPXJclG2bN
LejqZONMMLe4RrAVgOdsmDGJkDNo4ktDepnDcz/CdI1yU8O233u6gnLXywyYgqc/yc5E/zJWbYzw
XwiElsoLwMKGstctWR9bhEFiZvlsppyL6k/PNdaEdXbGSOrKm4iiWOqax8tR1zkcEdSr4n43uBhV
Ldh0K3hcj2C8zbC0GbD+EE6sBAb7Ji40WK9Ut1gClxTgrXzpcJc5twc2A50qcMn1+J60ihNE2wmE
GncZZcPRdyNQ56+KOGT0pzEZHrdkC92DQTlm9+12thh+nnQCfp0quAvtK6+daCd/Wr79yxEsSwTb
yr1FiektUFqoLNddEOFkYuwmBJJQpQC+gayhxxzA1N2Yheap+pSK8LcW2vFwyxuu3vMWGitau7cK
yvff0kLNOZ198uY7EZ5TrMUOvLUmPvRJBWOTF38LukGli2n3tEBlNk/HJID6WfrDlq6h5wHiRcpm
MZQXFWsRRyBR9vR3Zf8eoWFeB0gBmm0ex0tfPJLDgZOTzyVLqrtVRu0zixlDQy0ARtYqFYx6Ez03
hSOdFLM0XWl6V3Dfs96LqYZoXp2UKGlFibrdFKh7kibVkRzqH862jXrMhySuGzR2jHiDCe6LHWU7
7J5mO78F4mHrtgqqz+P7ZeqQ3V+6hAMVm6PrRdpI97xCP05azU8fDpr/04ceu/fGt4Vt3CuEnHvC
DIC2+JIZk3i3esIIf/aWUp5aoYb1WTUjZRiHLyhRdR3vvfEVjqbsJwfF3iFDGoyzkhpLcpLAOopz
pWf/kWlhD7BYdqIjtc73/lseziMjvSLi82xeiyZH7HUt9pj1t+eUTwoVAoNlS4g262e6W1jdcQBv
3SRYmvMu59xLXbe1imzHaVjKBREL4frAQWbgCneYSMHp/1pzcxtM6C4al3siVSTFKlHKRB8UL2q2
IXvh9RYwyo+p1SAKZeO/u+pmtcNzAxPJQEs9EICl4b/i61KP98HIPuI/fYCUDEJ5a4gYl3IUcC3o
bruBpJQmhYFri5wf3/nYwqg0+iJtuPtQvn3pnPLGw4SD7TZ5ABqSVXsvuwCzviKB8f22uIAPzqZ2
4UMj70u9ru3vw2qkoLBx20PowVyUuwUKJGvFZH9Y62xwzw4+spWireeX2LeVE3ksy1oKGA90hvHx
29Kpo88XscXAzbA2Nfe2PwnlBe/7YDcNUxHFV9+LIIsF62PGl+Y+lWB4F0/+80Va9WS4Ag6YL9Ty
4q4b8LlHd+bldFdhtrs0FVvl0hZxVzms61eDy2tqVzWmzN1Zer3thupS+qrl1gRroAcmn5NF7Tz3
uUITncKzI+T+Nqy9hKT2xTPpvoEgW5KnnmQ8F4R+v9L9ejY0UicFOWHVRvTA5ghXBaXWsPlHok8G
aNpak34ARsWETGQjn00tRX+U35sunfVfq6LPdoqtaOvXA230EgnSgs3SR6DW1SFhk+jP3EGEG5tH
qdzvGyzhtrEQotB0OGFsz9Oac5CpjoPZgT9dTPhbcpFMvvpYaQ9JtuMQWliwuUCNc7DZNJRy8CSp
0XLcqIolG+4DeZ5jTpqWYPQyeqdudN+zykWaOKS9+o7hud1Xf+XZA4UMG330kOHcCmgB/24gYcdR
pD3O8lm0ewCL1+iuHihZU1bp8kWIFUDP2R0nhC9al60+UFna1R79X9pJ/M2h5TmI8FYiXhrPBUn0
xVcLmrhhx+ujUVEG8C4WFVVBaXd36AR3vA2EHomQ2uUojb8DozbW8w928cHlkYGjViaXyhX1FkSM
uGOiXXMFjOJcn9AUr1zsm6JtDpilOM+J5/hTGE9kcl7q0YU+E6yFicaSFL87mV01ffaCmLNY6hjO
XbEWVT7t4sqwukNLm1nOckok3Y9PfVOpumHG+iMXsmYT1lb2WbP58uBfHLLrs6g71krI4eF8rjwP
SvEZnlVU6BtalDlzF81ZAsIiw8zZsZr6tdT7+xAb4Dn9hXm5V+K7HUnhCxrSaX1DL8xADaTq+AHU
wL6RBx9LOyEJCMvqEQi3Xx8tqvuWjeDMPjZnzu/YqKlCnkPRrUrNwcH/d1GvyJzopaLhpPtGe+nx
2oiun80CLFhC7/8IKSrxmQl43A51Lv8uz7LMFThVRgSRyol9ARjoRKQZ1i3BbyZo201DwYcHML/Q
xiuL3JOsUk7bE+oi+ZnR/ZZMYYiWACtw9v5y8OU8SBmDi/g/DE2fINAOGf42tCMsUua4zTePLrcp
zrIvygL8ZnZ8mFwC55dYL69cWOqTsi/AkWWNVvTBiUBOHQKipgAAOq20QZcR58qWMOWAcqHc14e0
H0A9gIizOup67gKTU6bxrgW07y+U8JhhU1iTySQhuJvYpZ8NAnDzokRq1gKazNS/AEagA6fDyaxz
TMZMaGHnK3JX6PaEDkcc/V6Y+y5wVUuf6ayC60FWQ4yBmV6cOm+iYo6dZEdFB8XAN6pRQESziuhQ
WGQbnYin48V/d4Rsc6C6h1g/TzZ7mTNf9ByyzLSlShGsRfrdU2zgGNMW8qHjsnmpFZGJ16edci1a
gqldI06nzhj8vhPVn0Kcf4oqNFzNhOq/AnTihwpz04D52vCJevuIEhmJWGJN2tyHIW8NL163I4Sr
GHSDiQLzUNkGAxwJYVkGQHVECb66t+/5M8d0lp1yeabuHOOTPDUspCHljV/dZSRGZ+vZ2+v1rQhE
QQH01u/NXKHduhFaBgldw+GNkFmih2epufWcaJGtPTIoDmKVtGBjxO/h+rWbXi+JhvJh6XGnTVK8
egTN0RbpeOHbwsWhSVsDLQdDJtwkx5GgPXLbgur+v4TVf8QGygBYPEps/Q3FYogFEuBziWKdvdUY
GAmNo7Jo+VDLitLM+SNzi1ap8jb7eyrgcvHlPgFkC0PGhPrn95nhfVDiZM0k6JGI8HoSrVzoowUr
QEKDrXOktffqBlSaUtPv8SjY2bhYEb5j3fXFC5rNUG95ndecCfgSULaP/5nUNftGFH1vT+gvtTnU
KluOkACQTFeRurEc5PVa6SGJ3yQeBo9PSjKBLL7MdmwqGB2LkLfYt9Mhv3QZqXAxtLllGvuAGAop
SAs24vEsEEd95wMhxWv7on5EvFaiz5GLLeMbVgtXuFN1ZpgIDUgVWiXj414zdsshK408jxvIJVXm
OnIax5fmsRIKM/OzjjDZrBxWKjDaLYgvFUkmS+xA0zp6TqOwDQXG/V1mknZevpZrmZtGorhl7inq
FL21rsHvm8hBjplM13zbGS71PHYyUgG//fZyO7GdQZ93vs1q3xrB+0X6doyv0S9HMfRK8VHkIJ3W
t7G+GBzkgFcYFmfcnX3O0XDpUMTnkVthQ1GH3WiTGNS6sRf+CuBN4KCeYswjteqQrO3Z+PrFU1Ns
/47bIziYCRsHKhoxCgaQTgjBPaVr2L25tWnZYoHm6Lr3Ng/p1gkROQBWI0+CivL2kmetnty4D/vp
J/H0Ca9tkbpGN15vJJIwoOLBEP6DZ3We0dWtgy/OfY3OlbyI1lA5H1k8Flz1adwLkiPiWpSmMTd7
TvUxQpX7p0SgAR24TGD5Xhv9jxtCJr8t4tTEG+JSgJfHfL2dx0lnE/9hjFG6OfzrztX1p7qvAheD
o03fUNd7v63H6K7pzmytatjpT3xRSjqAIDu5Jn4TWOpd3MB3mloCej0YSKFqs3YaAYaayhiS6Pza
B+E9cb+DUTyGDQXn3k7yo6AjTt+yCZ19VDVGbZ8R8J6JA6sFJmiWym/JmXI9aZxBTr1SFBRErVqP
XhMUoT9TQOJKUM7pBQ+q3avqDGyH0S4QRWAZa2vZAl3y2m0X126jAeAUrr7tw68bL4GSjLw6aV8B
1wPgPu7Oj7PAZ95SY5ZuqGuEDtY7JSZs+X7PQaMh4qebTPHeV9fXQADvDdwLYWIWUY+4haF1azid
0WdalEjq11nWPUcvV9bNuChQF8J/QSTeECQsYLjnTOkIjcmwWn5OYVOu4iF06cB50UdWgQCADpNZ
XJaLKDtTi/iy50TrQIRM2xpnhNGPWRpOKZeXPjIQhaZKQB3VkeIjtaBMF4LIoM0q/Yb3otF8xpcG
pQWkvAJ4xNzvhDA5o34XUdDhY7+/CSQQrfmld+nfJFotiv7SVOfVmA2c5TyW+qHvtRmWdBGy4QNE
5sLX7N/PYyx96y47LfsIxGZ6Uwydg9yXFzRYH7yzvXXmM0qay9d0xVaw5zMI45b5St6+igj4RBqW
fPt+pPdr0bB+rDSve4TJ4e8lt0vqfISmKzAnMVj84scyhZrdTmSNs/c9xURwYhqRweJ1/I7OosTW
0jZSEYCHkz0tkEe0b+oFkLYMPPYMEI5gCUGiUFCV62Z8hr006gGY3t/8rpELmo/Q2GoCYk+T8KfX
kdsKXAWPeVzo8quGuH1mI3G6rqI2dHATAtTf4QTNFpM3zwC+fKhlYaY20SBnrANC8LyW0jsQBZqB
RB9rTDqHymrMVIG3KXKW/Ljn77wGBdm3u44BeF9yLa0g5wzqv2YXR42ooGVm0+7ksVDSNTbYgQCB
rVoD4cIaOevOkOGCeyUB3xsPmHEeN1Xu2QHo5ynxZHimMi7Vtg7nQtNPUIzP1n9EFBmn4GZOjSh8
B81PEATcN4A1DXzHPefGjShv2fqhGgWI7PUQIRuGHBkFXSWaCz8rE1QGPtySErtT9n2F397dwpEm
pO81psOHyuGbpM70/oVE4RBQE2+DmcPnBQQwfKyKtVtnSf+wB3vYxNlXj/jNxRYWbU6asvdji3yP
h4qiM8MvEu8h02J15HB51m6FGs5kXfaCgUwxM444B+sAZ7jFKcNCMy12SoCcF645RaDPllwN65nB
/ABAik6P1PsFz/+F3UvQFw9N3gfDKJumRKNPM7MkbYIPvuF7tmYZN+0dkJ9nkAT6hDd2H/VMfnsD
3/X4VeVnWYZx05Lq/Zxy00x7311V9WqouOifVs/kGD6Qo9dQtDJAzsZav4e/L6CODJ0X9vIRcbq4
iWXjheRF4EVyd7LdRHGjLSJIgDOooqCOiZzfREd8bdcRQz8OCQoFQtkIU6FcMq1scDVCLsEZpsMJ
ri1m4qWN7MM2QnPTP0i2jydxyEmCcWXn50gv5f0mtlNpEE/njN3qHyL2IoQxk3LpKzQpHkbxAgIO
qtFFYwoZQ0P3FMIN3BJusKklKL+QtljpyWpPJY70QBegENTZ8dgQBwTsug5Cy9HGtJQWXu8acNqs
BwiM0pSetAJL6kZEWenZXYJ7PKH+73Fq0PqajlD+KqXCpVGFtFMXDRN6O8nQ2Fkhbn0o2CCIv3yD
9MDbHZtFwAPJV1rNc8VQ45atmZdGoh8BowM4987TyiSGZ+OnsmfZY28mhHMdqZq3FQXcRjffEDwk
mYiMFbN5WHyxJAkBpT4sFCIniqH3Md4NxbI1aCiMrKHzm/f9EejQWwBG3Eh3TpgACDGyfD0scMl+
m0dKJAO67s7aRpnQzOEF2ezC86uoFBwhnGwTDcm4A7EppFJnsR+Z6L3k4psv/XDIpntNyJpA023j
lDseLCbiteHB9S+OtMMp8XoV7Y6t0+UP3QJZtGrRJ38/5ABCLesvsj8iDs8pOBNTA2c0nVaTNJqH
4hMWT4HCG/I9QVwFDXQl2YkLWDVRxBH8rtn7MT4FgKFKHT5m8HB/aPBBSDnaffhRma4EelsZY5uR
hD31Ane74uevYeWOKUppZ/VJZXAxWsHmvwTFjGvHxu9pqUwneCmD5hVwuuqmENPDSRJMdc3d8uF2
Ufc+tijk5pIbYhJxcUsdn/ALFrjKPCsi9resltHiqTqm9C2lGyLPTu6xf/acXyJSV6X2tPbVjA0W
Gz0BIOQIRmJ8QeNlk3TbeO/yYlYP2YI50Rl03rMfpy6n8TyeMus34p7fLgPFTR/oJfjKXV1YEDx9
4XXvSRiREcmIRIw6xU4OPVXBDI3grlIsS2Oyv6XOv4J16zgftnqcubb26HfSKdTFKW3UAvoYCCJp
zAiEGgzHWFvUTUjD9zNjR3TnmZVq66oy1P4pCw44MGqwI7X6NegfGhTixp5UZc1QVbHdnyifzHDW
OfQh52X7gkX7H/pHrVwpxsu5VHRukgO6dNI68xb8mRkeKSvPFSeys3J/rs8rqatrQL97kIN7MWug
upU19THoxB9JXToqy2sxW8BzCxSKX7luk0xP4e9m4LVANfEqFHEmnOHsPvaVytDZdRwHNdTGVqiH
vWM0W9uyBKBIJyRL+exoWEpxPMSlGs/WbUHBnAujDW+pSUImS1R/e1a565nilIUfA752Q6CNQi+a
347W1p7sK9pat7u3wz67GjY36pZxfasLHuxIPwn//BGMHPlC4ARwfAUK3DIlQYA3btWGUzHbyzMO
ju7K13+LCg+WKw3G0M1aW8ACfAY4xXPgWu8Pj/2pHy9s633PfQoNyw/cOUXmRUz/pptIeWvbIFnl
Sx1xQDuuLsLtc0f/on+FQ0rmr2oUtOpWE4Ec3zt3ZfSrMebO55WXrnZFTKpExyVPpaHWKSPWG88w
KIIWzELpYWZvnVVxh8rebiysYr4bwFqg6gil3zyxR9NkCwqLBRw7r/SS1KeCb4oeqtnt0svJRZRx
X5JNwNaEj/vRC+LlsXpRDxEKWkGqV5PFqd8eLQAmL1zFEejUVj6pgOwwxuuCKBP+Af0cnGBh4GyD
WyaeMtXlMI4ci0dQ0lQaAE9xO38xINFRlSME/qGXRDJHG8kOtnSQ4dMY+1qITCilkt7ur4ua6EQR
GsTeFQLw0K4zlJodFK4iirjSqcXI3+5jOymI1dxw6Q2uJcEW61lwTqUrzn/byW8l2ilgfgeLIYtd
OogueEm+CIaOZy+vTFak5W3oqEUcvk3pgLyZCYfg9dRr6k8PN58lnVl1vu0SS4pYkmiDn+CTGVYX
GQ45hDAOon9KPs2sMHLfKNzHwjcCrbKt+9HALr3xLNFdpcGDa1AXTvtI8g7QIIO4A4HtQOqUakmF
v84laZ2Q/WgOt6eaIwgEKd2XZp0oxoQzTUF1uYX8HdWL3Jj9k20752cDoHaeA47xkIb6yA/Omhaw
0VTYSenQqThrfweOAxdfvSxq20h7MNdPsgrPhFtkAoJdNxpxwVu9vrhhLe0Fwu/ETUFahCUmtOtD
Y+0hbNp+7m7o/CNLUQwqXd/FxiISdYlbz0DYYnz+k8H1gaoyqqLHW5X0Zi9aANZpbFIpwhLnzyII
ldc5OLdn8igZ/lblbuO1LUGh8mVIbDfHK7aAxRPq70TP6Ytd1TUkEMdr+X0WQji8Xry09Gye8VKu
9kWU8rzAQof6oAaWGOaxNM8yYSy/mHsVqaDQyZvT4n35HcfoEJJSyLAGTyzyUVUKjcOyzTmlh3uF
tkbET0C4cu4EAdh0bh6eTQMdzVGSjMgsHFIXj44CLQGItJodnRdQf/7aOwiXwnoeTWNfROYrXdaK
Be/pRN5tyelEMfGzdVmYt11B75VQ8AG+9P/E7iBlb4gQgHta+m8Ia2gidWXa1huDrDvyG1Vv+T9B
4n9L8CtiaTjL8AkvCk/7lsA6uvATZkIHr/ArHcYMv9OR25vgsnkd2uLn6kMkfBCxSpGY6y/EoXhS
VKKJKb1t9374lDEq9kQWp3IH4Ez1nQYd4zcDlfORz13gwMia11SdctRJCqOXwh+Tmnqhyg359r5k
bqubnTq7laZtMUhXp6Le6jyuiq2JVvja75lc2nvCE0NKWobgm4UWwC3Ek1RIOqqHVNvQ93lqSncK
vit6EQRHp1hIKYMFlKuUUsQ4//uKHJTojSJmgOv0IHxkTDpNUMryCzl4Y/MLYNHQWxv0v5hsJ9Tw
l/L2RZrYwP7KywR1K9rXSv3cVyFGU2VgByA+t8lO3YVIdjnfCvmmmwUf7BReOw3MYDh4E4H9vEIq
ITlzNw9TCchM0k5gwDWKfPM53Q9IcrwLjnAswhDeBoeGQSK+ZvwK/1rZOg/xgbyYh1Rqexjd9Uwb
a6MU8pgLxjA/XBNlCWbKbgTxyO+lqr/689RMXeJfow+BOEU+2Fou32CbQYg5Lr9q9fUbKnXdTwcp
h7JogSXo1Bc5uRMNK/Xrr3aINGsQ0MlubbuWLM1cRjTZKGDFtXsTMbWcUwauXXdTabTmDjrtqhRV
X86Vw1KwmhcSR2jGyTDeMwdYyqpja2hhBDoWEYF2q9GJfyB4nrCkXj8mcyGav/9bih47SRzXkhBS
xnijBXLIP3H3grYPL46HGOaM70Ps66bLMVQatICEN8rH688SiaBkgvoAiMMnAmINcOrI2eqGk58p
K+Yasmo6ga1lmLm0AqVwDcx4Hri9HcHizIfx+BuP0QXVokDjIGqAcDZFr12jVQMKeyQOPZYo6xO7
sQRukzyj82WOQy/Pequa8+oMiylMB2bl4lHokeDGvT12LJEjKMMLQdQdhBNaADiequcLlgIxWQbw
Pm4mSntruNYmuBHXVzn4l/Nq96JHpRJ81Q16vPYjXrr7CNQIBVTnIqbLZbOQTaFXpVMmYICUUTQC
FTh6zseOnoMAxfG3QcO2kcu6MvYvURNyc6N+NnXcB/KxOCIsGrMQKJnzfweqeK+rpODJWwvRvoSx
7o5YOx91qWH8xtMu70fnZJVLgbonmWLz4xrF8zflkQp7tTBaRGhCoKoCy05j/maPBBl4bZE9+ag2
QtiI/KX5+10NHunlgDWQwr60NhPk0X+USb3wScLRFJlT45VRyyrYQXg9DyZpzNF5Ijce5gvVPwnN
iPaZl3V5JcFX+lpKQsHFOBSVgtIw6P1eAC/6Vguk/xuM8WjaUyzdL5T+3ci8EZiRaTzTHfGe6yCJ
HWRLpPt8N1XbweOQUFF54I4m/OZ+zqqm4k1AuE/zwLoRkcUPjT5yrNmbpxpLsq4M3PsuW3tILnwF
6IYHJ4xSq6qzre57ZYbAX8UiD/vIyj65qOdFmsHIUnU7nEfeypEZ+1BfwFk7kscSJ6UtMWLcVUDs
GwCM0SjQD11fSxJjcp3xUFSLPsgdMCIEVN0fTTdKPI/2g7fswuhJQgpQFHjSWq0FbCrWch+RD6u1
XhsdDmF4epQWeTZXcPZ3phKqNF6awCNogGA33rFmcNUTAYn5A539DtqnyI+xcIlZj7wQDsR5zJqK
MWWX4bPSwKVmrze7r5pm/qDvhtcA9cbyqKMaTHqvP6hsfz56XpvqcZ5VUlcod2ZTkQqV37nb7ggP
Snw4XxlZqQDfnvYf+ZlPREBQmBxMHJsUcX4+rM2LonN8h58jUPHpXdtM9NylFvms5oa8b0hp3TfL
xgUaNFPkWcZGfz+uPsBRHs0JJgnPmUGUNkE+NtVO27dM1Ut4RViaBeE5uWaLNiXPligk/zrj8NVG
1j5lLd+w+98hd8kI6X/2KKv9S/TBwaELSWTOTYpKttWaVRahrEeuuAYBAWQj08byRUF6HddGPyN8
8KPL6uzBq4NsgRGmwInYE4TLvwIcMI7dEVAbu2TiSmnVzieiOUve7dekbrPqBdLrnKyRFcnU35NS
Ud38w/n2untfjglIkHDqxBoxHuW8Ul3rDwwtZGMwbZbG8yCSfIWqk1y6PvBZXOAHVV7WjmZFl6DN
AZhkSnYZ/GoAt7zD19DzJ/DAmTmxlyauFepjl8fYHgNEDQisdgAa9uH8WBlqxxfX9liy0BTVa2/R
KL+1MF9/TYB3Y1v6hQHC+ARHqQOefEuPYSAEeAIz7GeoAehVQTG0qZZADWVk0Ppghx/FIKEOKohW
dt+OINF/hQqjecD5whMp4lESFy8WRE2qeuRSMdm30Kemw/diXGqx7jXpdUbJsMjv3wcQT38OCn2u
BW5k5sB8cl8ddT2DRbo/80R3CkhIDC+rybcxrfjc8GGYjWPXza+uqDDR2bp30Yv6LoM9icIcdTYa
xKJMVt/Cbu5Mut7pyQo7FL+1Tt6qyLOz2g9spS9chNCMAVV6B6RBw9HcPFFZQqh6UZrJ1ql4ikMp
0mE3SHecwRC8YUVwBin8OQWItHH+OMnefz/dbJFbYd70+J0YoQ60E7wOrDQvttcq1T++21rlKzaL
Es9MQT5Owqwa8m171CHfrqu5B+HFljFoLIdB/bNFbupycGloRecfVkhtoAgpz0ERFq5BTOM4QUMx
63IwalDEoC50dwbCGYrbNlmwZzMzO6IZ8PFVBP7+XwaQP7UqpDX8vzd4X0p2FGRjXGPTJPCsQxyA
ISP0bhGtwQS84TzcpxBpjhx1XFKEFT+ulHkTXu/Ny/5wVWhDpwl1GbC6I42JE3+Nn3oI7fHlNv/f
Bo8GBpaigMeBG7MFHcxeWVn6raa1EMqbSHDq+juHmBcXY/29YBCBTsiY8cuaTKlk+YtcmVlcJFOW
oYqgDEH3KJmGzMOm9Sa7FwpkrcZlpxFA7v9Np/LLlpKL5qbpUBfOId1Y5LInYtGkh2GU1BH19kt4
SrBWrv0O30nBOOOfmbm5wKohT37uTgZYVU6i1eqIuQJwUXX9pJP3+2oxT4UnTqmi9QFhD9gLn7so
Yz+Gn4qDVHhY9e6/y1hVsTE8LZr5PwqUi3mgOjun+MWGlls0m4+OZiq2pq3YfTZ/gWC7gBU37Wpf
MfWSoaA2rgb2N+u0SzgVZlFrTFW2+gLcG7vES5Ot2DRGMbU5rnPx/nBFlSfacavKS2yVP5c3CEFK
iGooSl9xWiVUFo7mcThCUdqEet7QFHYJZL0kNNohM28mt74JwKWlZasRYWmkFA5KkVsWYEI4pyJv
1wghfJomls7d/nwM44WYDZMR7dfdCxAAiyTzmm+j2ZO6sahLPwTX2InOS1jP9ARCPmn4VU/n0xtU
Y9DooX0R6J5Wo7Masic0E9nijt0+cXednODsJQeIY7wv32rYBa/wFDK2hMfFZr5Nf8JOI1ru//0/
x5IrWH9uyItE/nLC4lztOYvCs6EmULaJEOPc9wnPODay4xqz4aiNzjM2TPfN5I4SlBSkNycbVgHC
R2ooEazySV/fpdhRpyC8rnnAw86qaHtwPUhSJrOorD5EVjLv5va0QHbVuDXrPPjFXKkmesTdcQAv
irP7kuCvaJD4l0KUXmfSGEVgK4PERtFdGh5MpZgILwdnLiTdl+kunu7+qMe6N5vY7+nHQWbOSmhN
uRbL3tqBrIQDd8IaOqi/oFPxh3m4gj3bAdSkpzw/m1fzFQFXJNBEG58Ke4kGLCVVeFo4H0BfCywV
Liy7NVLqcijJc1UG70qS1uLs/Z5wDzms1mt3RPg3tbC20sPmrUTx7+j1FRI5oS8wVcl78i8K9I/a
PS397UaS6FGkVSvgGkpU8PmDJp/v/PBscV9LmN7TFd2UoiE7aYPWO0PMs/TQ7M4p1/eBLruIYnY9
LYsPQOPC6QwDQP7XZm5PxPCVp8gNc5KooJYURV3yCXo30DbcHn/pcQQCG4HFoXapZz0Df4cOhNag
kD/zOKOsTbx5fzioC+zJEfu5c00us6rQIMthHfeI2G/Kybb7dh2ZhUz14nrcZy5je7Gd2KaPE80T
PoRBFm/5sHWjTaDL/KS0FlZDClh4CthTAwBT6JNvYulwaHN5q7XBQ8RBUKe3pBePO9Nu5quIbmSc
GoMUdeksgRgE0CmVjD5PNYVYJMOsk2ffxL3xdfzUhbzdtCrf8Nu8kj2A3Wuk8HQmUIAeX4wuwPWZ
UASfj5tT5RG53d7n5b0aQRvox9kHNEJoRNYmsES93qFrOWa8Bg6NAg9DZkAy2dGibonOqtJk1uG6
PoSnTfyRnmXt4zmhIIHR5el8LCVE9Hz4f+5/2hBm6LK45qIHjgwVR3+ZOtKAXTppq0eamua3oy/n
3lNPRr7vAeFcdYTuShuZSSwWSTFePQ2abtVrqWr3xedX044nsbTis9m5ihSsldyWMrfV0+Jq49LK
4ELc/yIZOn5mOrjzjrIqkr+ueURB6XUtouVWL8t91m5yYEcNtY0sGprE+qewkIXcYWqBkmZGVjfY
bmQb9o/5u6im5DazZ9dWc1adL+QCoJXWAC6MaPvblS+rOkvdccxKaOjR/W0oqaGiJOfuFlCBtnxA
P5yGQebMJiDgYGK2ddKG+jZUhpPFFXqSWDQ9rQPkuC38tTU9cjh2/VZriiSArUzIrqKV3AMubzNv
NQILrUCExI7zwiodQT34YRFr7Sg/tpmIQj11qFQsfAcBVTyhqRjpdkHWQw4qsE8+B45zaneFu2yg
vT65jj8KmJwnhAIx4sVsLriVbFA2sB/7SsbyFf4BGUjyxJcclES4Ys3U9BQwsvt396ST/EShC13z
6YgyIgeKHlsrPnW0nTudXbzhetu4eriy/8Rcq/RgoL1RxGoUswX0tdIWdr3ccYB1r77QsATEDkKj
hnQXP2B+Q7iWzHgPf4OCG3Ta9Lb170X+c05JH2rHpwYFWm+WxxHbzxYKnXk7P1iZwKdL+RPVr4X0
p/yhGFbWWR/EVFhDXKwJm5ueDVAO9EQAp/7yWPf8zJkBUxMpMLFEhnZauzQzZwT3QF6gOPUaHVr9
VnF4W/oSIN+NQdr38/3CwGbAMHmyOGM67tlGTPXClbHR+3kknWDFCrtqbEcbPIcLuMJY2DFxYgmp
gnBZBPpvnrVaJ8zcl0R9f4J8qeRdvYTDEZW8Gw0iWPdZgQhkMidXRe3V53M76ibg5n8y8f3NhHDs
3z6cYkxUzEj2xxykLmMa5HP97LVnrR7llwvWs3PKGnkXZW7/Y+9yQtbmMonquqsKLn7DHMxGIACN
AA7mXp3d0HxhuKzRA0AFm3NHzkPIzQ4wyx4dcwqm1aEGQ0ZfbGbPCDUOGW6vCgM2o1zaq7htpd2m
1HCrUS77XGISCQU2cKF8dfN5WCKQmaoT9T3bQoBpDlhrzir7X96Jf6zCo3ke9juK24KvBBaADQ3i
hRqgdBWf2VeIS7NEIBJPOOMk2l0DQjlleJ6oQEywOtr6n06x2dME5l0ZTpjId7d+nxKeIEBMFjOe
jWwH7++XS1Q9glFixpsFo+H8Hm30V/ha0ZrZ/6hQp6RmEUWEK+ew2Har51vyVk661FtvZpI88kEg
LEx4/2Lm2up/1s7Axt4QOqbsPXlbOERji4cQzDH7sd2yZBS4uYm6HnkdfZIKF5piFU95o+eTRLLg
3Q5Lyl/Q2b2cajmQGK/ZIiHNPYP08+Go4pXRnQkuVjBesn92bQVolFSybOnz+7ob4iMQHHhFdJAC
h21etE8N+DLhIz8pkZLvXdpgJlcGKSYpi5zjIzG9GBQCcSja63ivRLVZAX+A7GmUCg9/YVPlJ2IB
m/o1hqBhL/kc6JdXBbUB7LbD1D3IMhWrkuK1JdecROL2Xze8YTZfWWy5lm44gFwwAJGfjBC3Rdl+
CgXXOQaoIiOi0rxA8KTvq77WqThFqaLFH1jeksZ0ysUV8z5mbA42qZSTLJ/q8aNG8B9reMJ2BE0O
slUjUWqEazc1c38PFcGP9sR8VDepaCSEzAbvFmsKpm3MHsk4H9+AS4Tjb7Fi9+E3neFueFwgKat3
ueisjGL3mTdztae3U9bVI9Jt3XeVrIlLj0FDjbQh4H9r1hCyKGgw7Gk9nxt7WuW5wGUcHrmqk/Sk
kdHFrrc6ipweSnjSu1/enPx8cJn82r/qQ3eby79ctDZZdfuKoJ+//cia5Dn5rSSFp+ht8yAi36NM
w/iuwy89twnMbz6eVwXshDqM6HIWcHrqieSWw01V9nC8Tk6n8we67MvmhPvv2WrNamlls6pLdVr2
uljUOk+ca/J3/PmxxoIbMskZ6ITQNiopqJOMx82BHOXGkLFqgFHAN3QK0vMJM5+jR/EfFd0tQlo6
y7g147SYrz5vqr5ugHdcpdfVnmiK9NdATf9S+hsXji/DYVIdLWGaVFUqe6922nRB7bpQ1rAHHi4O
/PV2Knrdu7VCZE3masyJbAl0EXfzbmOiVPpt3VkNB1jIRC7Wg4rDlw/ishFEmuNnaYfXDJSnhQYL
Fi8wyI7Yzu0unSezxdZc0B+hVi0g5QuA1Tp7kttfHi8XG0Ofu5ud4S0K1fZBzKfNRT7fdJ4vNeWm
8045MQqHX/ZzowuQpOkU/XfRTECFbeyn3ouJkk2yEpZ63mKYOVRlAaevGmrM6ksrPqzqhVF2d0TE
hdVFhkOm9KwVi8pyWxol2QZzmhtNo58MoMWWmbLLYyyVnP4Jnugi7p5mHqzJpyEUFBn7YCEtIG5x
SqYk/1vil4pk7c9uIS1zP3MhYPgv9MyrsV62DYuVb+jRdSV0Zao82BBPTsZHj8mhCqJcHGc7aDOT
LNxonlJkSYn9xc9DEl8lu5C/j/24DGxQfNF2cTRNecj5GXDixhEmcX/PDEts2xllf46gtjukbnq9
IhDa3HsTYGZUaLDBv7bkz4i4cNanSjaWY3YDX2G+9B9jU5BzpMKC7s+5KKNlstYjUSdKjKgL6J2l
OWDM1iVvyXx5wYf5OEecV0TUXv7fPBnkO4RjIIGBIWmfWEszAmwq3TtwJs0hKYqvEbDz7BAHQBc2
PG1sZnMCsD56mzZCs3vQhfkQ4sdyQOyDL3Aj9KgbxX1aB9oRs8iTbhTrMck6YKEudFJGLXq2dXlw
hDDj/iwU3GprNxW+Ddymdj/Vt4q6NtuM+IGdUbB8ujgxkkZVdMTYvr+zNbZzpB0ctmMehuSy50Sb
L9yBano67nG510UcGm9G6YQkRDuRam6Ua5gdvWJaD4L+1BLIBKHgA4NLFDnqEkB/pKJwyO7NbpKT
VWvRVFk5M7rHGCAfLbD0ORKo89aQngBo2jeR5Yl/YY0MK2RD2KvLrRqfeaptyxquhAL1zhmJmaYX
4RRiE3h7HgUFEypamIvfZ8EovSix4Za+RyRdz8l2/vQOw70Ix7e4BXWmcz5onV4qGyNkGRaMOaW0
uIwOxutc5Md1tOdynEIWAh6tZHfLAcb24d8457BGmI+uDnD+Z+Fa7XyrrtqAJ3ahKKK092x1qghZ
mB7Biodq4Caul2EqrR9zX7bYX3LpoRcyZKHWjGzI6HRSQc39X/4D1X9zWSucSHmwBv3qiSbe1cVY
oyy7Yk6pO6hNF1fnxMuDiM8TaEVNd1ZIVib9dGNBxcUMLelw7wpCeTPAp9dE6E2IjzzpJAylqZan
0FWat7Y1A7ccTTbiwlNxR/zzHzB2ZELlJUd02esixPHiVL7nsw9vxmkOzHGVtFA+QIZ8zA8H57Lt
66Bz1QK549qJUQnA1Tk48r9cTSOwu0cuaZafR+F9Ir+i8WLVH3Hx2j/Sm15XGoSwJen1TtYAnVfs
b6XAyddpKoX16Agh5dLMouk6HFiEDIfnmxCadP3ZZM6hS9tpAvwZmh3QwMQlGoPWOZ5ej3KD26PF
17+tdjVK5Q1WvlNIVR2FZZA8T1K4m1ujDwWFNxoPZM+Jg4mTwq6yPNPCMZHd5YRRasLLF5SSIIr7
vqIyX5CawGiLsc7c4wzRtMYptZqJsuUx6TFgCAmf4QbPrCvUgKBbi+EGbcE23HzHgiooXk5wg+tF
t3rHe8QvNp9Q3qWl5ipMD9C5rtlXgftQf1e7W+e1GQNlzhlYCPo/keEIFiKqYWu1duK63UMuOvLg
1mIK6aMAvLs5bz+o//qxyYcbu+xIoQw/97LPBMuBdvJgDUpC9oUGuQDFzOIXDmjLt7zY/ix0Pcym
l4nuByzYpMF+/H5kwiRMOpGz4pPmcyMIV4S7FGFw8mDiP55xMMToBkmGm+sThcITPKD0OyBvTl7V
6Ss8MjUQIgAuWjIESnJZ/odyNVqJujuzA1PTZJHhaqXAx0kTDwohBjsO9GT9KVvNY44RHb0Xzlye
CsJMOVzCIZq85U470H58czdBsJNErQ4PLC/WAL4zbyHb0o0JewRKU9TupN/GHXNSP940AuSV1AsI
4tFTz3FjCFc8/B3TkC2QbVJPAcf8gd2e2IW0aZNlAnaOKh2kuOew3RkEVhcuysSrqf5WbQzKbr8h
UC1UAO7xDZBb3GXwPWTZzlh8nAkHKrxrqSjj5u6vpTjRPKHYe+YUKKcIFqWfTZDnv0EHZRMUWIxG
dESmjSXWTBp/a0kHJgiQFymwDBWKDw0gbTLluwgKD9n/fEF0EM2dfI4spd6ryak0yDYeE8NLfaET
9CD1MMh21SmbwwvXYIl70bhpIaDSI5skj/WYsfdoQhTMYmwXPjzhAywlyx7c6vK4JGLPNQhtcXY+
Dq279fdEigYphPpLMmIAEglJiEq9figGXhqMyufR+b4QmyMtaQHOgF4+CCRDP6nwztEZYjnaMAUs
rv4AFffSUgoefwBxU/a5BZ94HWqaYZaO+utw4f2zppWmh97h7IfC3k0cR+f//UerlawvwrA1m6vh
qWw1pvnw9f8cRoophAUjRIcrfRZHP3HEDERUlY8l2jzI7+YAMqzXLOdQL7sMgW0H4/XyZUWS/aVX
2+fMAx4kugTWRsz9sDct+3bD0pUFtQbTSdgNQX7pbVqyvT+XozOHzchCKod9EMLPdoLKFiI4JF7t
kxKK8aSbhOh9TEGDDf01hl+odH3Ys/dWUE6hzprYyW5BLSBOnyQHohTNhyUJA9uy7Ptw87bAczis
Rj36pG5+sXckFV3j1mmh2S6kTNyeyQVJvUVj4468kgg9VwsWoY7SDRtHzHQ6Eyt5AS6Kr6wnaX+T
JihLpQaq7cUJhZAlSN/SYXCGfpKvu3jxdevewxg1ARtGBx8MXqGdXS43EIX39t6d8GEzD3rRwgsZ
CSWMgQRC6m4IBDsYNNmjY3OR61nB3K5HD7YzCcyoTFUdPBAsHqBwzfukQaSsTpgg/GzslBChianU
ZcqtTni0Dff8sJPovNpYsAzkRqHzlWtBOURPZXwGvHCk8b1525hDNzoQ9mgG/NoOsYyEvhCi85mp
shkGEEGLfyQVQPIY2VH4p857Gu7YKZSrFXYo0DJCUkE6+7Ojg+/r2CwgkDtJ0l6HHkguL7eyVecj
ldaJ2i008XImwoE6SuE+/ng3MCSa9psIescjd6Dg1VZwJqJQOKWfD00afXZBC+uJEPLAWkboPDdN
7Q4URKXrgGWNxfR9viwSrZIbnexAjbc3h3cC9Mm6jOgYgVYNCeI0ni2d9AuKLpmL5maQICqo4nKe
v6hj+YgYsGxhNDV133wuHXWA6P7qrTrNMeJDABD8eDJYznuGF5DyepxVlILAJTSDv09Oy3ZLlwGN
XS2/15p2fF1P9C3/FTys7Mx004GrcfB0u34f7e0XyhZcNwLJLVXEP1i04LzYRMb1znSKOIK3sP39
yhY2Qdrf44SiVL2AEoqZ4rdD519qVO8qzBMQXvv3DdA1MhKA0gAnnZBzymo/+4R4at5lPAjsvXZK
k1+eQ2V5yeSstSxJPc9dyamTdjGz10DaRHG3XDMyDREu/+Ga1GYblGeBuPckoqgOEukuyAtJtLzu
yWvvs512NVY/aLND+C9raYcfc1xCYrjXX0ImlxATyXG1O4miUbuXv8LmC1aA9wSffkafH4ACNjAX
YZAFEZ4fhACGxnJcSfgERnQtuF/SMsHVVkWWuN05YN7xU1Wp3xfk5AvoaoxuoIuRbNiVHcjRwmg6
qpkf5edxDRrRYlSXOYoLvqxPuho3zPJWluDii61mn663TKz/t/p9Zs0iosefA1aP2z7KOwiBZHYN
nDQN2NaPIpGZUbmj+EmVr0oT2mJfN9FOEq8jwsvP+WbYHyyV279mW56Jhf0DMG/1SQj2qsVv05/7
2RSzu/EKrgOETivVPOYuJc7HLf/aXzPcxxpc6WTiwoeIuEkPqodOnbrPjNzA1U7vWuRG1SPbiGbf
9HW+cRJTxNsHAmErooL73MfybYjZp6yrhvr1BxBQGnMxRsgb+VKFJ97E+xxCh2vzLi1zsvh6t5I2
74/kzeqsYyZFrHWs4MZRH0NXohEhT+42JH5qN3TFUQqwywJAOZNOedYyEB6g+0LLbiWUDluqmqJU
N0SOOdSN/Kwrjbz8r4FB8g2TZiFf+azfnGTp1m62f0mz/NuKGYXrdQI1I8BFNJ4bgGodMk+saVT1
QJ8Ltn89C0zzBVXcEPgyg2CAr+IAbeYy+bjj94Mx3hQA4Vu9ZD4T7yHkQc8GZa2t52e6s4V1Qkc2
y1TKRRMeALC28/iK1JkoL2inlXVFi9PEz82VD39JMBXw3KBNUsFh/SGFX8E9nFspnYKWdH/FrpWv
gbwabvZogJ1zGo8X3duggm493n6Iky+qtDvOysnvM79hHXu28pvzMQjSkE1rS+bQ+Gggur1Guw2C
L7BqfL//KlikQ6yqYcBffI3KtO3Ot+rvXU0MJrP/rra1y5prF8nj8CpBnjU6C6lSlo5oteHYisCC
MJMZ3QBYT5zIM6YkFEnpayDYAsVfIZEelD0V7DIgXZImhkcg+8wphXWC9NYY7G4PDDNe17Lm268V
usZDpJF/319pVnai7Brfrvdvg5qrb19HRdzzsRywZYIIs4GUvvXsSEpuSJs/R1Sny0LWiYs6vtbW
AN+D2kF91EB7p8n8rB2PtliuGxJrFwfiNkYimbkF+TshFsWnO+Fwq9WXH7hcDaJiE9L6SkICmnby
GnlJ67dujKEw+hTzzef0iE/EXsgdLSYI7lGbD0l0R5IoDVUcGcr1iUxw9EEvLdlCKiH4NxEkHQCe
POUIkebtDQDMZC8EK/RJA8CrLjNP6uBHH+oICwf67JyprHNMVA6DD3VLmdD33dyNQ1XZrJ7wcG1z
h5x6r0vPRSMMtrZa0z38Qo/bpwatWGIh+r8mp6UUsgIN5aZKT+1Vikyf6gyd3gKw0BoPWfOPJM/v
sjBWvKI9F5Dap/KXCp0WYk4XePTAXohT5ttyX6bZtwZlbgIla7UIq609r2S3KNxI6PN58L5LFXfo
MUdCcExEap6rEIs6TsnRgt7G/6PUAsjVVnUTqD/4xf9f3t3QI66v27aaD4NkIwsZHvFuN79TEI4E
dstsUF+73CHAR72z5arQPL0zODECLKMko9jueBRMOJTy44t3TbTyEcrVQ4sXhGm24TxN/Pu2TZlv
Qm+Vv4FuinPZo+9Rm0C/S8q3Iwd949DUMOU+GCFTjuVZyEUksfoz8X9vrZiCo9Or9LEevAnMQYvN
R+ncQQwU9AliJdpX7mrKWURK9wpVbljM4Cs38jG35TZOB7pR10v6IhCONt0WH2e2BsUGSQR35NGk
M1DXvMVO4Oyagt+v3LH+s68q9AveKFpTAs6Q473y18WvAtYrLZCmnb+DfyBN7B8Amw83qWj1RopC
O+IZ67GeIC+MU9jPg3+THozFjAPImmMku3qGyz8dxYSMRv+G5i1LSyesl26NqXpCde9FuB5nJ+pn
25ZlzoWipHKHxhZhCRrImNXpQzt0Wdy2sbPDavCn3iF8aU/v0ApwZMX2wIrLbkJTbUNgf+TTFOFa
mmseu6k7xXHViWM/FscI/fq9fCmyZgmf/c84gtCdlXckr8gM2o6JuX1Xdj62d/23VFHHBzCY1wd7
jhB0akfXHQe3lY2pFyX/F4Tfh+5as23pYwxo+daC2kxLzBFypKLoVkhjztNeznI8WUQjL12xv0mi
p8vpLNzcGwfxXv6AG6RXYGYdoIJGKpMN05x20zurPm5HjnFYF/TTAnI0YQqBIca+yE7d7H7/ceoz
El7vQ2uR93jfqh/57He+P2sTgfgZhK9oQe3pv6vUdwGhXh5Pbdxba0rEKV+bisOgBA75/ssTxkCR
4/0FlQUYT4+/azBd5JFUt53Sb5+y6KTSvkJpGSDewXW16JmgvobUJPZrTwvx7pv59lBXgOUmgXJZ
Sns9MgoQ/yvWyivYpNHZ3lmJrGnbUb+53R1Xdo8XvYit9atai9mm1RQl4zzhLrz8bjWPwIABrDcd
QvsvwrXtS7QZXy7bjQ3tVcULrkWZupuH3SwRr3GzvKE5/2TcuY0Ekrw7JiZSvb8ZnOW18UwEbidc
IQYqijX0TMpU1gxsjqw+C6wruvmqSDkgaxe0E0l9ukrMfLTbI7N6E2zgwSIjlxIFE9kh8Iuhmlnn
eOxR7o8c1zW/ed3JczEZj/zU75A9HNl610oNoPBPRo+UHfNAmXjzUezDeB7xMY7b7TJoAZgxoR89
TFiJ8g16cKGptoxj+JWGtkKW04+OwIwfU3W/He6rrL6cVM/zCsHbZ1sIkcMs8z6qQyb3jUCUto06
+52LHLxVxF207HzKAZOZbUJtQKobwZ/IhmUD7y8DX+hGpRDiuJOFgnCi9AMMZDq7nkQWV8ryHCFC
8k0GPSzDZmvQd82ewY7YzE74DPOK82bIqUFgKhK/AbM0qNJmmgEitafjaNXbZeaxKHWcTgw0l28B
AdtuNPvzyy81aJGgCl6+LC9ztBzH2xe+zAfUUnMeO8yGLdaPxlIf2QXnqk2XYREW8fInJ6huB+bT
5imFI7tkzo5MGcEHOs+PHUdJT5wRV6rLdUmhp6ybstukPQcA7HvBqT8UAdW6fgPee09ssvfDQtNj
ZqibQ3C52h0KuTAAEeKTuTsWe7i0f4wox5D6xaT/rcO8VA4djrXfik2IfrFlloDvHIw8UW863AXT
yWRnsStAluujJWhAQXGXMJIzy8sjRuPLfFU/ka4CaXMy9JLC445sBPUIZaUG0mUoSwKtmGRWicW9
0VF7x0vbUc/OLxjc25xRCfhVHOHi5fIANeDiWwSiM0yfIDoegO+39eJOEUKopkDA/iN4Ek6IqkzP
wutenqrm7XacTkPCbAL3FE+ZuBTk1DUOifUx/vlR17otwoH/iEm4oEUxNOJOrUMZ2kyB1MERpzlw
MF5psdQPjBN3JqeqCZ3ZkHADIl5ib4QmLEo+QSZ3XIAcjZTVN1jBxuSLkUq+E55QUPzV43AOeJMC
Wga4Jo931+nzbdFEzPsW/c7pxUhR7nv6oMsA+YWgRYfKQv3KkjwsQVHhypdNvCQgfZlqFMGcPVsG
vOgDWvmgKt6mI+qRhxgdsXBvVlHQY2gNN81bwNGESWqhp7TNkIQ0mXdGSAZSGuA5SKiLUWvJ8yFL
KgfL/I9ws78L3RZAHwL5t8lZMPoaXSflrViV8oSVFlq4pPlWB6cUxhnoehZxDKJ/+8KnlUEiSTSk
tXgjypNju5/QpXtzVJasLSKGVxZAZMnNgsiafSjju2hBuzkfkELP0lRBNpKmJndP26BwObwoj0EB
IzR5CgJdxfteZ92Vhxphs0MrMcy1mDSibthLC7MKTCubDAWOAfUKaH2mSZer4MqsYkoEonT3INEe
+2vDmNz56ZPih9GAtvL8iYZfvf1J4Z5yiot2T5QlDwfOFKGT3swT4z6+JPFLrWulxMA0RoO1DYaM
ySfo52RkReMtmbp+Uam07MilNpK6spkDKQAdyVgfr4UsASmq/HwRwNdtoAi5NVwadmyQ1tL3YY/h
4ud0RGFT6DL0N11CENnyhkxCjgs44RSIjHit9+LjB2TuWkfvMqAg1t6pMDvwN0sb8SFvJVo7uOJ6
T175R7pcQrhPbV/CYRXpaJV+Z6P/9LN8drxeCXxINGMfJK876mH1tj/1cPYmwRFi2g6p/tnHfvsF
PhTpHxQTG6ckWZ3a7lGqp/rRMshcQdB68RIlgoeFRwlSuLMvrD0qHYi6WLnB6wLUPeH+/cSC/qFa
cH8TFaKpheJrys17sZimFFYKnInEUnmZdssBzP7bvxnpwkM9l/OZrP3RnzuUgCU/6JVALWqLh1e7
DQV8wbJbkpsniPUlXfkvIPlJMfxmh0nYptbDZFqGtODMeWTnb4BLwyDt1YrF49iAX5AgY+6zqkqf
NYLkyOxDsh+PJW8LsFLOt0x6g8mNFdETfGktwWOBmtP75L/9tM6niRWYFmQCKpebRtTjeqU0puIJ
kEIjq8HfxmKT562cjJ4f9PpZ7gzkc2dzemcPO5UkYjex2mp9uG3fRq+U0ViPGhgoGHaDwoc5RyRv
3ggvStOnlgVgaUoZDICXkCydrt+w2wu/hnFaJBf1jF5liBi6Je0fx1ol7FsSd2afH21A8lAHZGdC
shCNLgpZZ+YA3ULImi06diSn+oUkMsgA/jloMxYWXWeICmuauTgqb2n7dvNPgHNTVnwere8iCFSl
b48h+ML6+1AKicVeuIaqtb96ojLWL5I0MckP1d68b46ycA3M33lEoSlI4Tm8i2xRX45MINqYmCHl
YnBSeYx5lU30zjNgXdTkwFSEpPbc4DSB/dyz06Xa3MxTJEVD6b+BiN5oVaymXdCrh7qOHf+cdDTB
tuiheGDBBLRzVwNsh2UtCN6Gc7fDSmz1hrEoLhCtDPjz1J1X1jwHP04l9VQWyqUgesG8BV+JzzlT
csNwWsMfQC7X/Z4WvyvWAtjgFSnBU8sIDiv4X/VmPG+apET4asDpI0omzByN2dk7UfF8ksloRajh
TOyZ342oHmqPDQoTAqnwuFKJbT4ONJQSHTC6S5DXqkdZgr6OBw1aJ+D+WhdxtL0y3UIhPEA0PEI0
6K5VKeSYV+mw+oq+XJlxRSzdGl5ODwT5/gphHgwA0YcgQ6Q1kYtN/M325Vw8t1TCQnHnIo0Huf3S
UKF6ilocvHjG23mXBNNZHrl66ZM0Qg8UrgicEZI26qg7AGZpq1Q3lrx4ikGsckxi3+2Ueu/unbHo
/xRYBYGRlVwtW2YpRBKgBClz8s9YDvlx9hYnXdnZM9YDPqunmp1NH4AW84C8MqC5Bkjsvxfy96EF
yQSja0it31PNRX/xJRKME8Pg8qZldkp4rM2/U8itjWazZfhCSEGVhJxFYLyLy1GI146uypBHCjON
7U0sQ8Jit/dVmORP5vkPuW9oQnML+DT4Mb2B4ovtSoG9TiWotN4s1/QVThcls0SGx56rRwzr/aOT
lHyoCR3vCqzLHj3u3eM/m3Tx/blOdP6dn5rTYNDVZeFpeBjq+Y1d+FYgc32Z7RhWDOpfE0t7ROei
ZbSeXtJ4FBu8JQF6+PgErJuL1WTDyBOxwVJWYAsoJ22lFjNH9jr2NnRX30yarSU8BkwOnJy8CKBR
B5H8jpwJ+H9eh8uryvmfVGJ2dDkGjtxhZ4/hV3sADGLNuPbDizV46acq2+tLnAfqoC3v84JjsKqF
tI6PRPdVd71jI+l+XE7x6azOhq3hQrvVQCshRoMKa0unYa/EwfIO2G5tdw3yrzzQ7TlMCZXFaVrD
rMbKLibxkY3LaQzkUY7tJGTLKnOub879iBOLnVM82nIHt2csznwU+vjrbFCklq6IhX5hbX+4LAye
IOK7BCgaMWaMrko95eALzX3FX16jtbYFEFMD/LtST7p8mJjmHHZSgMjr4KLcbGsnjcaJzgCJPQ8o
bbRLVMCXbwC3IU1i7ZNNNJgkIyoM7me+J0SiX+xbuK5pjr2ks+YYh1TqbWUqj6IPn67xb7vp5V2k
2/qmt8kw8Bve/yiRW20dIDUxIFSHxzqDGcrEy5AvGvUNTt1axg1hwO9CsgULcQnt1u/bExpY9Hn8
3vDcF4jwzN17ECGj0bmQrY+6KGULEZd46jznXjl+nU4+GjyeyNa/kOWjtZBTmL/3ywLnkVALgY+f
OM9o0uIP0mpLI/hL68vi+rwO2Z0JGpnCadKUtAPI3vSy2PBKjKZd5VoypqEYtkqko3LVQkxLZ8iD
2VJxKI8eneCDyiYRbexx0J4ZONR9pWBIRpGthVtAjzm5yXW37aXPMAFl8FLNCGLfQlVJFktNOf68
+LFgm0/hypFS+zHpy5Qbohpje5t6OKzj/drJcpkMFavqbLGgGxlDvcBam+lti2l5MfN7jdF94czF
Wx6WRLn2JZijbDoV4r3AyXWNGN8iEdoL897oSFlcmIHoxTrJthC8Qae79vF5LNWiscPYiTB+T1C+
Uve2p9GdFFlIHXcmNigoi4Vcf0yO5OPDxARcurq49BJOLO4xyIwX0iXnMbZogt0U1Y/8kcF/pH9D
u/MX6hRYIYwEBRqndiRF3xfUBsqYQg0weS8D7ReJQOJSfQKBxSZUhBCMLF0aszzIqaI3K3lxGaIn
JFMVCUDL4EX8bVm+e18doQqEqsaZjA2ZgqNrmKey+C6ChtCeIJ9aqfKbA3tUIfzUEcQP0HqaGbKq
NYL1WsFNSt3bUzOyB9bTKdt66lzV8Rs60pQOLgsXTGYst5bcd83FeRJaWiMz3hiXrYdFdS49p+vo
ThxZsqcqry0e85hN/uaetoNWFe0hBXHEyNQDC4rjZ0CfQMIVleLsFD2iK4pJnDRyf/apd937lfBp
zc/xRkCZ/nJpm6bbiqcy0M5vcO+pBfoe4xgil/ob+k9/7cyMB8S1ftEK8ALihFYzi/Nv3P0gSpNy
L38CIZ7E3rmY2um5iih5kuoVyt3ygprDIllkPzE8j4OZnWDy5HHWfpQle4QRqX4Olflq7quCnD12
rJUFDMMKxs3gVWsvmPmTqZTtCsrFaFyqwwAtivKOH7GLYJSIAFe+Sz/VZVUj7HSUR6cRgQftQe4U
RIWTva3XOPjhoBtHrafl1rau76AuYV0uhYtkKRadkEK5bkWhDPsMww9gGqSJr58UGRCzjZBZMYsH
H2T37zMGxpNMNi3PBMqlBaQ3SLp/scNJyYNPMSUFNSi+uFjxG9TAja8cOjzQqtI3tPFZtnmcDRoG
Pf1T+OkdGhHn6MfxrO17xzPcNfjjG+12BbCqVun/kgCQlXSB9TZkCLhopzS953NvUZgji84+3hJh
ui3+mGluz16iyr/SxKEGrNADZeBWTisV9hMaq8TViLV40xGBMO5K3KMcDZDbodwXzFCw5MQHM0NY
xHa593A78BlClCkb7FmR8M1v17kAoqqCUMQhAFiDSDWaBumqQQY8EjsqFG8RnsRnXVV/blTTu0Fp
sX/tr27FWVeOw7/5XYcyLO5YVCIoSf1BOse27JfA1Hs7EPVIc9t9g+sGqTkSzoZe2feH4E9f7wP7
RxBHKm/tGJNfSRjp1Wyi68wqWr+bw9FUeEQR+o4IzCJFxYPUroLgLj18MlKPDr30fJpw49CYltMZ
27wC/feYfqarAECiYzrRZhxr0YiuvjpHgvMigxzZgDTYJSKMjkD97SRIcoUxFJVPdfikjkx4F3vh
PLaiA/0G2uNixgNYfzcqekvMTTFdWn/VdZ8SwKAjCaOASUJsfpoD6HXuZDiwDPhT7wyeosyctBZI
piKfxiLli+MY+rcsK9fgciGIaNKOg9LZaYussn3oFs/YfonAJN+gSs7+BmKenIBSPtIUr5WhxZW8
/24TV+jUfCtFBG7/Lj5B7IDvLUxJNWhNa/w+mv4Mru5yaW1rk5sObrEb493D3AhHfBKHUQAK4Fc4
p4w121T88Odd9LJVEB4OgrCjq2E8oq50LtX2r+ugLCXaZgTbGwzhbykNzO6nLNSHFXeCDbD8Oc03
ClqQ9NO1qHUgAU2jd+jdb2jNrMkyoBEBTMFfmmhqvsR/R1qmwYU33ozxnhwknyrIzNeHwNce4cn6
8/8l4thDjF25KUTAW30Q5LrZCBM5oEk0e3PNFQppRDqGK31/E2I1WyGiHULtFL/QVuWk9HIrnPYA
VwfcvGLieoHaSdF9KDV6GARoOnwRqa+Xoo9qLHn+tGuk5iRCVH7Dglme2X+yobw/0UUgyCklHOOZ
PdFeVxzZ7TH4Z/RkcD/NPFclWTy3sSZWQpXlQ91PMCwl0kNjAnkfrzalUBa7RQ4HGjUlG8TP3ZEh
kJ9KkBRAB+ds63mti+ry5je7tRKB4YWoTY288hFxSxEX5jdkOPGQ5S0q1un/glEddQZtWDaItpjh
Z25e91igsf/FkjXpAci3DTahcBYr8Yo5x2o6BYCDJcCmf4W/OPc5OPnm5kGt8y1WEQ0tJxZI7Tfy
vnUJpKxUP8Q5InD+wC8K8ZdwG8U3BfivhH7K2+JBHZHZkNnaDdammhY6z14I/v/sBQnB1d8YMJL8
m708FWL3YeHUDbPXzLNaetGk9CK17hEo0HtwclybNQSqzdk0HGCwcsWcJ2pBVMxkHOIXdm9oFIda
zudMqyWxBRJShrtdn1frBtDZGisl0QdFKJoqyo3f4fLi92W7PdiVU1yZmuhJO2WI98zw9BYAbd/2
J/lj5WTH+h3F1+fWbd+qz2qlUWl3Oo9eIqF2J2iQq1J1aTHFWsVE1/KUz1p6YHO/58/5pal2Gcp0
Tsnc1KqAcsoCpqRsAV5ZEWJZKiRvskEBvlXY7pV6u1iTdlkGzhKqLwwupJrEJPtx/y36wVrs/Fnj
j9jq1JzBYBlbuKU4x7F/8LkYnuuCde7Zxg9v1b3//YDTkjfDxjUKoHUA43CmiLIfnUrQEj4rlHom
2YITkw4ozjMIt6r0jYtYuGPoWEiMwdTM3N9uQNUpnuQtYiiKqq9azpIudLkE2FCwUY3X/Kooslb3
PGh8qSahwNOkucIn/KIM/n2u2IFDPC5umMst/qjAAUeZaKU/jIlPG/cqmDJZwLeJh29NWNHfRFkw
0BdJusn1CpOV3gVkuX9zGlanccY9dhEPVISXst23hFVGxrc8Xmk8ot/AHZRtC4c0aaC8tYmR7U1V
5Y67xqeXaWxgWCca7KOBS4s4ZqitaeNOmVdCLZvfoUNT1jBy0sUrJf5FmqAdXkvIFGhVD5RVCY5h
iJT03YkEoI0m4LeKtU0mdBske08zecfn+ALY+PTBRJrc9fBcEy6f3b4aUAg/AAyjyTvyb3k1wdw0
KkwN8padynQ9/n9dMR0X5AZb51WtT4GPVfVJ4av6vwas0XDESgfQOv2B8Kwk3wauTReukWBU7Fys
SaHUldglJAsARbTnMgE7w5zUnhs15/Qc0DxAg0panHJ8v52IrRJgfCJoYWRNXOIvhvl8dublZJ4O
LEqSo5F1ukv6v8tx0h+XE6iWWJq40TWiPY9NXQ8x4hPsjvb1DnNAad2UhI52MDSR8S1vJRi63NBt
m6XehA0q9RLe5Xu2uukYLM/kGhO9syFcdqowCSa2vivuSXOTPZ47IxR5mJamQxkAr6IaWZpROngS
TZvZ4i6InUZlICuKYJ3YPynyqmqc7/ZuxFvGtE/NT4oby5fT/MMY05rv18ir5MSw35WCyOAmkedz
WpFxaVPz+PlXMooLJel47UXVpgcFj3abrFsCpgrOrNZ99B2KYpaZ2IX053YpvIKsLMjmMbjbHrLw
sU46waaYMNQ2Ive6vA9nysDwIIyibcf+3GoOem5BvP501Y3SDfAk+XxUSYvDYqlBZGgdklSMlvUj
a/mTGstnc6Sh+PvaadAodbDWplSz+zgvVs3+KwQBxE/1qs9uHy0pHOQRZD8OI15hkRKAYbUCuOCh
iVY1jipddQqNAsSJp7BYaNK4Fxhk7d5Ilhj+6MEtcKK9Do1/kQOe1zR+pKoc3bvY2NEQeUgUbijw
KwOtcXve4OpCZnTnhVGHu0oVe4S31PVGPK+q8VeQEVNglwRVM45xLbQYnmXu5sL0cHPBjT2jQUJW
WFwkpYNoWBQoUH9JokMsYy10fOo1/fDh/usBEOjyHqinv5RuxNh5y3pFhjyQiCubUdJFHywN6SZW
Q0cLGljO62+vsWNtx6sEAdMqLh7Xrscv2qB1cJctTWyGPOwGo4jNODeygkbSYtaWTK7Uc8OzDPWv
YIFrWhmynf5DgJp+l72ektq7nRsbCTRmJsLw55SDnEErZD9YYHZ4JRB+ec+vUaaWdyFqUJh2B9X4
QTUo9yTZZJEn5GcpazMVeBJMhX6ohkp4C9fna983wrProIJjUZ8ylUHQ+4Xn/3rnttuqslOQVriY
SZKksMwQJ028t/UnRuh786WkeEEhK5F7urjVRnbblSkAYxvE0/jkHPNlbwfmiAUgXZ38l31B+TtC
eA328CtXIwWbz0u9bf3vhtaqi00nDcvGGyZugMn0Z+44iTMilfbpJNgA1SFGj3/puHpqw+5ghefJ
6yFfDTnf2xYqMw8LwBfhfGl9XgSravoF1FyuOKynUsK+aosZ+AVvo1NIT47HCK1DmpyWtSL44a+s
bNyDf6dgKReo+w/HZSq+LEZkuMryq8ydhQPFvUcCAgVEBipmpsnlRohHWsnwAx6S5wmBW7iKB3JD
7H9n4LZNgk/c6R8xfoiK8vkMPQ2lmtxqPTBbX/rV1SK6FkOtnoJ6Z3rYUC+dnvT+0gGc6VxZTK1M
NQ7Cy+RdC++ir+blmVIaajFukFIvg8nqqsAIp8+1tYcI2/f8aZtAaTiXPFeXcindXRWZ02QSAIQg
xhUiGuay6aljmqENxhnRG/CopjDXUUMBNgsyqHDWXFj1hgywkM3JnEbVdaiN+D7HFwqyj1AZHnN4
gndMcyH0EY8kUnPm3wuM9TyJ0ZW0R1K6lUTUk0GQ1DguBZo09mCNRNA5HXD7HwrL1MfzS+r+2b7G
ttco9hQMq8BdTH7JNthQOdXsiBBTVvcHoipZiFKhgmN4X1XWGBqS/2oQSmp2Hzrm+bzlL2rdRWEW
idaO+Be9zNlJ++gDgCp7AkYuA8E/YCzTZTbvrD3sNrQr+TA0wkypeJ5ONBFeAu+h3OzjCXfgCr/X
yqL2BNjmN76+R31W/Xbw0LNe8vnT7odLS2Hg/MDWL66op/qYUqq+nLyVcZtcHB19XRWh1nqRKmq/
lAshFHvtGUaUrKOH5abEv9+9YdsMCB+vnHQSTABax+9RzM/6c0hWkAkj9dBWPFiQ8i5N6RAyBD6h
a0o4CCF44C8WbvGgiyGKWcDnQMewIUJLvkFNgL+hkdX6wEFGu0nBjiQqGJTTmvXRcrilskdg2EOu
PrcGSQE8xH87zXngUJnTpSDqTknTunQmDvdCZgCMnKNQgmOhXBLe0HVcotduprK+66uksdes+PKx
6LQef0+SebLpcwa8eDUAy1xo19VtjRslQ9qc0kOLND3FXkL7pk77Hc0vLjwMUvlfmoFB/DXMPxFc
3iuxb0Wii6FVRdq70W3I2/RgpuE6wPKg14CMPo8lqmHxs7gNH28eh5ev3zO3LLNJ+R+5dHwOZyup
jyfiDgfXGJHYzHhXiASWj6e3I3sSwTo2OR6BuXS9YZw1tqiEEszxPKo2u97eoD9tf8bMo16wcAuH
Gg6o0fmsLfkdR/mZb5wzVAZYkz0/gzo4XyI76N6WmLwFJKSYBsUFtW9ejlAL8yliZpdiDF6ACam2
Fv+qHKhnsRpjjWCT0f3cKmFJl8r6SCmvlShW/X9PhDz/4uKWk+1/Y5ahCykXM928tykN+gaEilMD
QhQt5OCz38WP/N2q1TXPAx0haxnMzdrJfCA3z4cmWUN+BChhT55+q9nsQLZ98vkG597dP4zfMzrx
yiAWOT6Y4bUFyxJ/indMbxaWe7tNWsDBDvcE59l2MilhgMWV66He0PyrU9S2qKr1kJ8fp9GJP2Xw
iXkn0h4P//jR1M6qHDpbhbF6IWuCJ9HMehvjaFzUwxC6PU0GkXx4A+E7Li9vQjNhv4I/8TyiL7iT
oEZ3TQihziTcrj4ZJ7ge3fP3c871HNEFnv/pUVf5GlZNTI2JvmNzr2p/4FTXuZ7AfFanVzP9qLrU
EPWTZn4SZiclREuERCCr9sYzhc6mDzMDtAR3PtrPHPPez3waw5pbfh9szR+fFBqn10bLs3M1w4uf
dV/TJ4zrSbJMWsTYPh8dvcn0jCDmyMQ9Cywtg8c+xP8ur2m+ku8slEbQclJUdPlJr3bj4yoxonIX
OlVC5B+livk42IlcGiFlNOTeL06j6FNEehyLCyuv7x8DvnkiEGdqGMmeuIjWeHH5R3c+3KKvxRVo
9SgCIAGHhN5W/lqY0OvPo7cfrUpw+evt/KJLtYIBBIkPj45qjX0Y7C42FiQWSyaEcibCFLVXb8gx
DAmC9SS9ShLKfxw1U6Zhuohw1Va3VsJw/+36CDZwUVt+gd3VU3vKH0XrMA+5i8zzBls2pT/4ffp6
+U4m1TET4Dbg8jkVK1GkiiMjwoIipJBaBZZx7SzXYTTRNXSACNVeZLhLtDJlkklp/u9qSGk0VBo5
GTta+jHSS/sSO92+vXHK5vtcjo6Ye4IR83YI+1oOek+YQNuhnve9m+WIlakMGMC4vFCQwyJEf6gB
gr31hQJjrqmJYrx1hvHOTcuBrBuoQrf6IniL7VVtm04ZiemfT4azVqWilmVOGC7v8L01Un1fd4TB
xBwZrJfdjqSkhhqRfMGd4W0huWvqGMA5MJiq5tP8r6agOkERGCM61+9Ty2Xftt/26rt2x0WYsfCv
pflEuGF6xohqWHIkrOimfJGWsKJJbmTFQkNRSA0hA2aIx59RYYilN+auAh9jiXSti4juhFVgvmPO
Y4VSLUT7PoTKFQSd155SMcPDK3pD2LDsuyL8Rasl5vo/iR2yUtuvV11cuybQcwxIE/fd9tL37trB
v+Mm85rSgcOkGt0Z8eWt+26Ofu3Znh4JqJ1nmdxh2qhTt7Qt9+AIKSLF/p0hop29QA5KkM3ZyczX
ifXoJsTqJJQmTOKg7HNx1EtJ7nWRr+Kf9DT6ZksjVbNipkKzQACkQbtOnaIafRYXXqaUlUoKJ/vT
KceRJb6++L+CUghnSz1NVRQPK3wHoUZbs94L1E6956umyrY7MxFURgI4fccMXZTyr2stYqxh+vge
9JKpErZyfnLhyKinmpAotd5DFD0UE6o3dsPAY5SzXw4T+QUaUAjOwn3MDemHJUpNzxW6xlMu0DvJ
Zo23Bb7kpBiJjeJXhEgMxiBR/7lSrTCi79WHXZtOt3yVXoXXK9mJupyddV6ykUcu4evvYYWqmUqw
8/off0AybO9RUs9xD6bM0oFlWvF8/+ReAMD/q+rtJpYrrceI4nZC/qGJk/wN42Sh74vY3rLRP6dp
gZRmZJA500pDHCGJzztS+kUEq5KWtZ8GOchyluSwnAnhL3wfiaW0Op2Ul96Zt9JddTTmaa8rZK//
+TUbG9ra/OTeEAkxxikFDkmJTMT8TJfMX+XvKCjyvPMi1Ta5GGnp3N+v2kMQ1VSn90KYIE75usQF
8vbr32RNZiZG/a0QEAN/VEG79RulIgoUoPtD+D0AzG0XtE0XoxLu3WIo4+XlrVtkeDI940pdcwjf
RtqzfJIF5Sfg0bzTF+s/Jt8qNTmBBXTAGLt7Z9W5qUxmDTTSbVronXgV9dmGLuU3cnmnRSn2lUMu
bSpNLYIXeeMt6IW/3MEQkzMvHuBJy3hNgh+zYU30Usk9qZfWwtz0pabRSVglJ8hvTDhGEm+xi3dg
Db5tA3BTrioQSyhgFDaoJQSMG4JQ4UCIUu5FPWNcCjZBnnVp9DAWg9JU78yM35DfkU2mCbcb63wW
SFJ7I2Ei3Ba4od4Ei2XV8MrKmqTpQR2sE6ZE79d0B6Ah0CnynmPRTC3uLdYGcbyWNYnX0jZJ+lOQ
b8BtL8COjQugZvdtYONczsn6x31B1O6jLlVOSMicgYIaLFfQwgABDQf7GVgIN36P/K6Wd2ePBF5P
7j1GEoZ3maa7E3tRAHiduIqIatpQwCBXks1xEXDl1udRaDaggyIm/R3f+/GLEZbPkeopW2W/D+R+
zBH/zOsdLEF+UzNCwZZr1CJ55lbdPgdKpkXhanTbFbmrPrarzDvsxHzwQ/IFvDlNpAszStaaguHv
JEw3CqZdwh41j3fYVHqQDD2hy6H/hIairwUWzDLranudbKlzL7INBYNLDusWNK86L0lNWisAPq4K
wcsyrw5ddMPL6+4AaGnwPHyDmQm20/XvT8+zyC5Mn99wzKUeQpvvC5hnSJfC9hMxNatJaG/DfM1X
W2gOv4Eq/1J34s51oVBUwW5drfiYBQshWRpsXeEPktwzJoJNkA0/xIMSL9KXaf0KIU7myYShxkaZ
YStcHPq+6U8QI6QlvJNQ/QE3PT/Y88nT3k13f8yjZp/VQt+tQEiuEDzNjgSAPHrB8fSMXbK8AjYb
QZsJlzh3zkOt6Hrw1RNArIkR6ecrmNOeVcX8U8ILvGnaZY3ABxkXL6s7Dt9/5jWulU55jquNB2Jo
78hncqjllAyNzkbEt/CCLuqhzUtcPPkWLFyHiVgpuujPW0SNMbnNCl2ZzaC4dLGx11N1KBnKGluB
+6CgyHSand5WhLSElH3nR/kG0cuRfLIFB9ckvYfL+VGHVpweNPlzcnxK3QzJSOQTlQ7KPaDXqQhE
w4dG1jLSu+LAKfIkyVzW1l/olPXPrWJ7RggNuGl05P5b5DPNBfjnAyZjq43NugWYJ1ulBoQIwNRn
aYMgLgnaUkyIcNUD2ZgoUBfwKwox3SCB20Rp/Iguk8GaCjKWSPgCDR4hSRLdpDwmM1BWjH6NJak2
tEsHRwjkGcvN9C5fgU4yRurV84Ev0vIAHO0BS5N3eAsFyzIQyJJGxk/AToOLvyAUUzlqR+ud1eLf
McU+s38GxPgcsOdK1KHmixtKlgCa3/0YQhi+ZCTIcm+hh9UgvX3oxru6Zfsm5OW2kly1c5YZq5fs
9CMQOb63NG53R2GInPvZa00G1gxm99046djetvVXEtQe4NHG91K3SysMrAwnpJkGKV2/K3HKsyoF
Zdk5Gttvhy6cYAtzh/cyzycvxY1AYfHcV9uTNZB20OSyR/YVeBdg1TVYXXaYWvP/l4kdcbQmxAtA
9syt25byNE9CRAXROKxUSTVfFuUGLnU3QSvNiQNjz8yYuBPKXqBKuz3kXMCbs8K6YK/974Lsz/lA
pwjCe3G2/007wba/C2xk5OCuz3iYBLT0TuALbBY3x3Faar1yQ7l9t4JnvZB6EAk4wQR6I+uNCSTC
AcdwojE7d7dVBo/SX+GRkZajneDwWiehCRrOjo4giHmzvi9L0XVuGlFWUPPBKuZo/tyr/jksLD9k
UM1hhoxFzG75Y+0NdwGZ9lawIZl1iQnlBSgNgFSeI9LV4im7DPeQeiHHS5T7Bpvbbd6L1aU0gOD0
Z6fglXO/7cchHXruWvbyLwYFNrXYsIf2zhRAWBq/ZV9FsOxsGfA0dNyLp8i3TY6+R/Yk37bS2L1X
XKjOwn7KOSjUkD4LxYIKc0viWfpx3HE4nS4IqGg3ZpgLhTG5OMFLrfMoeG4To7okHw3pI8rYsh9S
WZ2ftEYu33pPjc7tVU4udTlSSq4BnjESpa6/04et1x/zNeKBhby2bALAvzKZDLK1SQnZn1amHsm+
fdTajxYJfimYMD2PHsbiJStcewVY/QHASrofFbaGJKIzYmKoveeq8p7JyaiKYDYSd1D/5j6A09n6
CcGrd1T5NWtjotNm88g3tlA8r5rW3rwTKUTQXDZDPoEJtslAtZpKEwyTylRGGBuA7fuKZmgpwrF6
QwVvYsTxvgC0KBAyA5SfWGeTj5mMDcCuCKX0ihWsNmXGPmy6Z5JtK3mSxYHP3hcX7g/W4zCbNWwA
AvorYOX4uIp1tiXpx1+rB9UGf6o6pM5tx76LUolAFA2jxkk2RXG+DRFwxZaj0AmQruCe6i9HZLeH
8lB8ndZHEsCfC4yjARxtSlhmF5X3M+hcoWls2Eiop+bTpKh9a5jTSGD7UvHYHzw8eVCeR384TYsu
tnWlVueJhYZ3Le54D1hSFHLzAYD5YL5OpYO2Gy55Fj92mB4jEQj2bwGzfcCWXouZi4WrkktL+d9E
3tkbHed/4aH/VYAsElCL0Njr4kkNbk6ggyWgCYWdghSWgladbqv+eCBUBrVfFATRHh6ItHEdvnUd
Plwq7Wxa+cL2geuSjJAeH/pQQmzptFUW9O7xrltP0+lYxoaLFpWBquUuHipGu2S3Ifav+XvOw0nK
UGHEbsq6aWoMVEKvFHAEen3nyBZ7LdlqEsEUSqubwd++OGylIBBJD/jtSHwJsUI3i4R+7PsdN+YR
9Qh9d+jn5G7Y5MIucwfjfJ5yx3yjY4RAvLUISL7F/P42e6sv7yMr6Lx3t5mfPEHfiJLWyXxYdfcX
Ol/KvkSDYC0R8XOiti2jEysbChktEV3NZ+Di9IiahAuQpviLvYY26EqNg1M2fpkQod3vMLXL09q6
M2p79mhY61zX96HxDjMEUEVxRljK4l6T7+0qC1PA3GHlHNSjgIXs008/M92xBD6VuEKae9zqzKyl
lVHWU8oprtzhiGnmVdh08jP3hgnT9ieFHlO67k1d/Fz6/hQN0K7I7p2TzVgJ2qXOrqb2l18VyUWs
SkorWpOyL3EC/Nz3wZ3vHv/litR0CdJfwdDSXRpJQqTR+CSyMjzWFFVFXoaAkl+skJ86nr3jtDrS
AcQh79CLisyiPaIP3uWhOGUlkTcZgbMQDL7FFKVfnbM2+HxAGniUjOE57IkGDqT4q4r5Khnc9O/H
oO2tz6jyhzK7cPAJ4ToB/X3cj0mhemILh0ZTk5Qz7qYTKELLOLfIoOe6UogbfXAdQnpvXhSQDhOC
aC7GV5alY4jc/klPxXbl9PIx1P66QbRCt+zskcCTiQ0yn2Zpd02eFPe8bmdBeG1nXBZmZ8KPB6B1
a67ehyrkRwG8ia6RM5Lris1As91RDdlZj11mc63pGqMiYI71grlsXsV0ym3lcZ2DCxhjNzSa08ee
w7cZisX0gaYLdFenVHpqoNUjGPYW65+TcptnucUTw4Fi+AcL66elw2ghwGpQyFJ+HJnB/7aowEzz
GOyU6B93SjP80Jd6MrGr5IKX4yI2cJxrfCBbplxjhhnwxL8Xo6871t6cjW3/0KcO/hVInBViUTDF
zmF5Q+GEq5n7SikvzNCtscaCwDPWuGF7L2U/XVYQ+j3OHpuEXs875UXOW6Sj4tCxPo/DpvbTF4YZ
E4+GIDpiVERUQm6DOQ+t9Ms5KqIe224/txnct0isCQQzD16kUTbdDoqJC6AGV/+ntnPbAcRTr30J
4CpgRofu2QADBVoXpLl57+imlghDpUJaNsfok5y64IhVvJYtDdgGTRsB465BUaJWM69XIIaBwrIW
63ImwKXA8hqf5Bgz9c3+1bDkQwJPH0jFbU5xyH5kG+xHF3rlEkuUVubM51DYuJq+1sux4B7lnl1E
sDJkkBT9hxuM4NX13tkj+BwBAXYKiGTYgga3Ji1KUeXebInBO0qVfDcUroNAd1bF96ec0hhycn7N
6lQFelYaIrCsaFljocC7WGrooTGzZTqC0j9XbjMk0OlguHwUGD+0dWqM8Y7P12jiESwLed4XaPsx
FKBIcFqZssFWO5uNLMhw4kfj10pLk6UxAMeemHgnhxoyTSywunLPDWfDCoIZU/oid6ngkz2HzHHM
dg6GlI9W+TnGuFc/QflvH3g9rvS5c5WrwZY6/XZiuypC4SB6PhrNiVawnDDOJGEFEKqWoc4gnV9h
5E/gDPpO7fYiJkDzgeKUdO+ebQ+sLsrmo03Y+D9YG8tBuG0Jupe+AI6hPsuP24Ai3uJovtAt7S4D
GKHzRqJv2WhjSvvXDVcp3lEfCggZ1hGjIHZK6SOIpEJiCga8Nz+ufYEX4QhKUAUvEOjzTit4bhNZ
IqqvGgBwfkzZi3XhhaBc5rvs9Y5JcAAnLc/BBy0yCrvOvRCdz0DD/Lt/U/Oh6sf2toB3qIByVaqi
VJFgnpFmNCleCBdQDfJ3Z/94QjIRijChjSfezznZu3VukfuGmEQEpigOXW5un8jSw3kd5jXtAaKh
bTwlqMxtFx8kpPavC6EVW9r9ofSeVW8Q+bNuURq80iXdt90VGxMAL/FSMzGVf+cr6XBKRX6Xt2Gu
RpwgaJ4fSLCUK09mqcqhNqzVAeLl57XLP+cPoiR0r+xwdSI2nUraLE6JQx4dsCwQQbWRRaTDGetd
B0b+/FDbGFfdiodwMBUJTXH2KUYAKoDkVbowx6R4pPLIMCXWun+97XEGnuq+UQvDPq3MTfkIbJrf
O2p340wsSpAw50OoxTP0UC2/1hH79B5MDuGsCe3Uv7CGoIweQMm56nmVZ+EcpMjVyUoOdFhOnJ4F
UG/rBA3MonkX1di1XIUELkXG7uE4EoGk/faUzEgWrgI3dz3Qvdo+enO2iLfdwdUJyB/5mXLqH/4c
/oB2WGNMC9DXjHX2omaD/iIpziYe0eo/PTLUyH1mb1k9Qh1veWskt/fgS0mQFOR018qFJLeZ60XV
as1BykQXvdo6XOf2xA92kKOa5/IQFsDr4YLztdiIVzitJrsS5YTjrSBjVDefJkOd76cnYGGZg4ql
KqqfcsqLnEEGW7tNJdfK6N1Xk3Ct3Swh8pe2RVohFEPHMdVZNFog9cNDG/WPen35mfkEiL7Hr1dY
wL6H86AGuPwQSDt9+xM696NA/s79oBzOoxyYOV+UMMe+aI5K2g4mTUgV+yjoOlG+zTfMwC9f383o
Xpn4u07Gj8VeCgJiMTdBeSR0nq3HzZfwLlEIKKdMz7w8DKwq6Kl/onVBgUxJUxwUqmboo1nyLlOq
z0mmirTZvc8nB7In0I94V9KEydE0tVSWN/rc/otWs2L/gHvHNG/fKmh3tQgqVsMRRArWomOkTi3r
YckEs/Dq86jkN9rIVG4f83pGxXlI1gOwW24XchdGKIQTJ2l//eCWytjzw1MIYUtDxW4Zh0BRm2gV
7gvv0uNe3L+NiolHboZJ3p8sPMVgyDDx3GCMSsY82cN1AxD06AB9anvfTeHtME9QLaq2dOYAOPpi
OWddtUpkTlivO1XcP9bwD5AfjkGHdsRjX0eBdg1Snh+Uj4hAz9+kha0peoudyaD2JE83kC9Ff2fD
pzdMlm8XaSCEasM42AQAGsE1cZRGdcY4f6aY8hPZhBXs+zLE95tkDGjsvIAEqdCfKdqe28PgzuO7
aR+PA7+PnylRsLgkoOd7pbidBwYGUNGP+9NXeFheOHLOiyPDnMC6HsNFb68I6Vo8Ibs0rEoGN3CY
XaULMQfeC8HDwqPOiid1JIK6eGzzrc5/EQQnVJi12STOGChVEoboLlVEW86y8TymEVglwemRYZDB
L9gi3wmGwzPYMjUacVLs9Y1ANrCNsQLS8eGvGNxwtRqxZjWJJy/JCCqyE3zlVuW8vKrmxHIpsKOr
gx4Y7CuwnvlJlFWrv+efIvfF3AX6swOA1fOL8fk2GPtGTItTHCmrKsUaD3Yc1aYiwDNXEeiioNc+
AQ+ARBnBsI6758vzQTy2XkgbHUvBFoE+oT2ToXNAhfPMIMhUhgza3Zj1vQPh+GdTGZEPsN9JIgDU
ZKxqbBumb7vwVVMc5ZxJ3PdWrdUSVo6lHPvYItNE8AQ4bOfXfr6QSbyhAXtkcONH54Ie/ksp/CBc
dDTn77afM6TxoE/66rd3a1Nq7uOi+mJatqVNoNmgHBCYHOeBLKR8uJP46DzYMFnOcBPBuTb3nQQC
e+R7IJW20qsQSq3PMdWxigun3eSLyvUHRfP0ber3o/WP0iEQVQ7Vwm5Ym4d+2VQ3pT/BhDM3uWxd
QdxLssQYANcaaZFu4fGnEC3OHxJhT9xGLBdY7XyYIDvz5VCaG30LBZhs7lHlf42WEGLuLJavIl5t
Pb/Vt6de/NunagjYTxDgCssW5Ir8j5w75xx9oeladN+TFg/9xWUtyRexH7YjCcmt/L5CNQpmnW1A
SeZq2uGQOWiS4uArXZUBBPLUElMi4Ypg6emFK4SJzU0aigpOSextNTJflwgAvJ/WvIq1EuBC+rA1
7s39YgCQ+SPVRJ3gTl+0Dry6FAk8q2SAm/r1jdr6epQImbC8G6egrPoN8XHvsmfIyuWTLkSw6Chi
iZhq6WXJ956gusREdoUExGhOo+og865liZY0DObmJV7KXJ+zH9rGkrnkvXrY4ZOTbfEB4m7LQD3O
fBWf09sN7GC72xe1bggQNB+v79aqyTt+7x0w/vu4BrgcyfefX1zHfGLlcCZtcI4DjftKhaXgB0GH
poAVJ0cudnyTdhoSaWiA48dI2JeCrUVcpb3u5FnU+BMin/jglsaI11LcXYuoU7fT2s1N0lbATg1t
37IKWzj6GTrRcFTLHqCJYvwv9UoGEp/EeCEOM2SlMEyI4kzt86c+4G3OjWCidzJtqQZ5empcbcZ8
Qq6jWKj6FBmsQlZ5icUy8llrDvUIaLx1h1pd2bv5VGQyVsmtzTarz7eC4PsmvvQEA7joxzKbHCNK
qz7b2tJ54entirGTgtf5XjiS96IZFeso4r01CQF0wgoXfzZka8schS/kYcAY36Nipt1IvOyjoJiF
OIIcWYEwys5xcu964W64IIFqTRzF07Oh1/FjfIsdPCekIsbNwa4+bzABsXHs3YUTiZmoULWgl4V/
hU6JKPPfESpxl1VJa4BqHoDCTPG3la+KVJ8phd4kYk3IZd6zfQJZ6iPTOb65plfOnYkcQ4n9dgAN
lQcFlrpWrqhShETuLlhQ0fx32rd7xBoEdWrAlo0KolynzXr2CSm3E+n5QVwOn2klXupcTSXzzSL7
tyT7Qtn8dWmaSyhTuItd2UHk4FtuLlcVjjm3WVedFK4Kt3l7XeI8kqMlECvBJv8w7SIIG3hCZIqe
pcWlrVBQQuwx5DdGhvUhnDhZNyuBiTPaQ2bRJOhNxfuLo/8Ya4Qe1aa4wqcpThcVaIH5wgN+JQRB
drevNZCjpNukhqj1/eqxDulevzqZPerjljGX8RayG5iXzLB5vg57y+fz39HLSnLQmOwWbxI0sJld
0JqKMJJemKhMfOjE5KSY869JLwaho2sIIfiAskqv3GP4dqH+3iTKfr4l5Q1kTnrwciAs+8BCawIO
p33ewUf5d498Xxe5TQHwvYZYyT/XAZrfxSP+NDPciIpLxLQa4pesoaHG0fb+OhHvjHhTRmeImUL1
W3J+8GSV+wfNdj2tnbl6ERNON+yDNI7OuJqwHs/NaNLj/dQdbUBZturG57UG6XweolfMrc/bLqoS
YYmL2IdvXKpq2Ihm7KF/6yu07Zw5hdqSkI0VvsWGva69G9p5dfXDHOEfPsBn6OVvmhD5/PR5saYI
VpJthD1lq6TiScsKfOOA3UuzpE4gJ26sHvJt4aE0D+q0JtFGDUOVMoVxi8zWB8PlvPjjs1bqQdjM
g9K/Gvrjz8Lt760pHx58DrbW4oN6JEJZxSri7lDJtUk6LRvuP+DbIVd4R8E0UsyCuuT09dzT9nP+
lYxhz3nV07jVdi7QYIuDVoUl5KoCv7fFZyVddqSkYjB+1L5LhkiKYRdkyftinMHTzPk0kMx35cuJ
7lypI3LiH35ElvAXOlWd+fr6DjwaJoLps0d4R1OcHq3LAkpthyw2Ycqg+ZCqULIa6I45qj8hZpck
f5O2hCr1i7ded2EcPkD9yTFE837wu4WJynLkmmrLQUqnA1dZABIwmDfHK9HyvlaSY+bgreqrYjaL
N6v6rhwTPptSwtjSxrQtfE+zzZzErXM+Mpkkya0MnW+mSXX9nopfoT3mVR66R6SRK3qAcyT/erJu
Jhbc3mLYDl0NDCZL+k5ZstqKx8sLh0JfgS2yvvGopdvpvGBD5N2M6QktlWrnHBo574uhHg1tQeGC
0NlweS8JL9NTrge+isBNzdBhFdDzhf0MmkgqRG/CSoaTbtOMK8BkId8U4GaVNULKzCr3NJKEFqih
f7HENwCqmMUUz4eq73Tq/4SCrSGvMdXJG8PtLpMlfs4nVm1aLTm3Dl6u7X45HvziZYT/EQU58Y4R
dbooecZJMPztDzSjltHbTQ+q8AOU28EYZHMR6hjHLPD+xD29jJZSXg5vK4lpF9DCD6eedeMQEgpg
BlhTnZpv1BmJvg9WXTesyqfKUhuZGqGW05/gcoeNEe+YPMPkY5kVnv6I43oUBwt7b0nADq5VMC04
v/16Tub1a31ah1wYBPLrHjvU2qxvaoZWEfsVxHfXruD5oJZ7K+dU95OXwsxY60x7oREvuCXQD5gN
W6eGF6wqQil/B0zyUNqmKGhDJA5yqfcZ3uS6Erj/kx6DiPpPEypgdtVGBW+4UE+kTiMp9Me8ChX7
Xf87+DdKmhUT6kJPT5FFN4MkVZqgVBPHKpNSME4tVEjofar0MrUsppWOR2d6VEaUUw/e9VtbOZ3M
8JZHSO1E97ymgaVo8MT0fPZaQEBi/0BAnzkuKK5rI/gr8lDy43QGPMPe6tCcybJUzRTr0dnaZjwX
m760cOQHCqAvJ5+zIEVfuLmykT/DPVxvsXdhbY9B/vyDEYJCQjrinGDyVPnkQ0FSEV0nUHEi+Hzk
wLd0jjRitywpQmcNEV1qKyHbAO20RtrZsAXNE9UIzavNyXeKvPkXr1u/FPsinyOdq5GVVObLkQZ/
Ypshf2yM9f6gqFzlnw66g4JaVbkqn+V0tww5zfq8u4eMm2G8SM9Zmz28DxrsWgKoJ53v7RIB6oAg
FGbBXF9cT7Ut4w4bAWBGdr7oSZJVVsd2+i7H6IVpr6CdezaXV0x4b63tAWXHNSwd1kTeiQ+UNOlS
MHzIoNXzb1rftwLigyxfnr6B8inLFS+sBd9eQTbDmoXucJ3+7lF9mMSIi0m5x8GwdGJCqftBwHiD
EpOwMm+F3bH9kSaJFAnSWnVJArVTSeRhVpkImqUJiD3elWBqa96YsmsegelOsd3BG9fn3NoWu4Tb
X5nUR/7xswv+2PT858RYkNxt1UCMIt2cgDIl/ckMvtpfrM8NSBRV2v/K8RmY8EsNExJ++6JfwDHK
6Xzxa+SlCSZRXG4CI+VSQIzhcYcfTh8goBKJ9A29O+mm4EjgNtfoRc7l7QKJchFIf/0dcclgMWWN
xPdDxocPeJdh4yMQwSpRl+hJwRGmq937qb0hVa7PhZtz6aZRjTYdGc1Agm0E0WJZBzszM6j8i8bQ
WLK4fTC70nb0OEWRlBlMITha5wbiCRidJuyxoRKP8bjDFY8HPONQbO8RphXxg+KPsqlDbjrl2Qnb
pv3MMG+FjvocuLUas+DVXHIkjNbrqeWStUcq08kTCJ2WN7u5TtiGlY6ngtWoyd1TRVUlyPlVJ+HE
l3MoTNL2DNLYAimtsLqIsM+TZwZ1Cb/z5qCrLf27K36o2MzL5Ay06EB4HuOZ7wbrBA4iOP6WruVf
YvPOfPnggCBzyUAimLdV919a27FxdGSTXRyOdav8eWo3Ai8IgjJA3S1H14utEYS054T+2xwjxlfF
13AVHsONDn3eIXRywLAje/9L75zAg/KBAVozT965vBGhukbG9qTwFAYR0xMlTVlALEoSqVb4s1Tg
/baZfSwfnnsvPkqeU4qrc6XHA88DVAMDaRMCRf/0fAvUgSXJ3pGRNamOjahNe5j09uIwlHRjYMnJ
7gqLC+eyezja/FYz0Ce1KhLvSLSkTl0qPj6IwTSMniA28gblLaxKSlJGN6cHQj4lf/NB56MlRxr7
V5aCNa7+QYDPPmSVlm4IJAk+eg5D/5HGY+CuYT3UQ1KyG+4nsv/9hL8RzoeBS5Fd98cspqEt1obH
aLtteKX2wUEJ0kBZhfo6WN9KqFAAzPzuPJ1P5X3wqLhExgFFysMPK576iGiXuEL2henw4YQNt/uK
NfcPRRHQpI4iwC4hC7I0C+cKQsgx0qKXp1j8Q5XiXLgZfJhX6Ph3eTxG0123rGsupbehyEAMdNJy
csaUH0IYPhbsNNYSDcVBz5k1K4BdQ9smVQVwWOG6fS0i5KoNrjAYEm/5X7jvaJFF4NymeFrXyTCy
G1pLruiqA4ZAUHfue+EF/o1X4+o42AkrSJ6SrtzypFHbglRckRRbedk5HTkGl0YGjIkESmOSXY3d
HVyp8jbntDY6c7SGebyteXdA1MZZ75Fsug0jd3njwUF3n0f1zPZyCkL4lhHCUl9qBo+9XSdobhLq
bx+3bCk61DbS18gqGlJR5CuPdjOXYlw/B3aOABOdvM3QEmSwS7RsX5oj6PpjKp9XQ1pJlk1Bnodq
pR3/oiLB1wfSEohD9tnRy81SNxd8crmnLS5Z92FUDsUP2r9Aa9xMlRiyYBI1yi45BXj3Htp8mnxc
am3RitzCh8PO7IosJ981e7Y3ck5Y6nGJGc0LdLrld774Q75RecA+pCJNADphuOhCi0G9cMX9tp0S
jMQ7i2oAvvAo17j3D9EUyUu858sZUy3nAAEVVlptnOA55OZ4p5dC4W0NdpfQ238tv7jcyuurg1lk
QxZetenbjVlPGlkCClCsZHNFk3CdGpvSN0eoSTjJYBPvIt0RfMQ8CixASuoAsXYMfs9VWYEKgv2U
kA2GI28Ln+0MYaeE+zvn/4Gxi+NvXqLmYtc+3FjI64IH10QUIVhq6kxfNNX/Ji4VsekYiZl6lLC5
imPhnzI/ouxhJSZHSO3gk9tIwmzMRbwB1BMVhefAh3RSUf1BqGDj57pdZEkV0YZt4DEHjUXFk/ga
HenKdpnPoyQVoY2B3FBNh3wWf2Y0QszKq8i3Yoer4AeyTdBX0pbx6leJePDDZFwiqJ8I4MzvjwS5
DbrqYKykHMioIL+o0MCnxL5oVv2OgrJrQotumcngkTzzM4IXIz5aPenmFCe+ohnmK3g8A8U8CWDU
/BzIyNuZm+2eBfI5hsZvfrEI0SzTAEuruBT2lddrLHHSO4mGbUubr+6R72/Ei+puTRVSpvnCDkhr
oWcwSTagFEh8PH4R+KPYm4kDlo8cUBcUAx82DR65z2SyCGRJIVxDDEj9MNK/ePtZmOFtR++p8mq2
xNmwNnJJxCJjlgLjcBL4kwTx+H2OwygtfQ+a4H4+q6eWQx0pfyHLmFYpexEObB+oTXZ4lFtbitxl
bBv0pNj6m8tL37VP5kKvGdTzI4Grxh6FQWN8fTL9M3KMJocsX0y/maDLxbgX2jH+N35aAAGj7Tl9
ko17IINLHlpdP5WdnIgDVZKSt9pK9L3ORXC0KsbBtCy2GzqMzoga6akX3WCMJaxMUzihSCR025hI
cCA1orRukZk8K6+TC9HvkZAcEKq4CDKr9gmQTx9dADv+xWSvzRRB1ildCdzeJbvs6P5N7dgHsDK7
W/58bYeD6ZSKTdPWbUNjYdPEkkC+PwSNFoEt27MFIsgl/OWpHr6ihs0khaLygaf2CBB42DHqn48K
VeSH86WFfsnB0L2QHCXyKybf8Fd2yGG9ovOTrCzWeVa7SqWVl+YOD/qkILs0Cz0NZPZjah/RJCxe
yyQ6rifZkULDcFhzwvGt5alAthCeggaWLtIs0xYTR6TP2SfFkYtdy7kwa5B7FlxfDSgKFAITeRLv
GDS/Nhee1g5CzlRlduM6L1bDmNiQ6eOO84itWQO5qIk1RstueNmzjpIJg+AXgPG7xyy8lgrE54cX
9zOnILaTwMTO6XEub70bFgfMiBVez5CvV0jP7Njlz2VyEzuuvOhbV4kl4JaTMe9XCZMcRLZzT80L
XLUIBbRmrb+ce2yOyWQ70wdYqXspuulnv1lwuK0CXEQ0/di9M61GIWmuM0HiSyyMUvSVPZf6mWrM
Txw2vei83f+PuoC0ynF0X/t/fuPxVG0Crn0RLIMs5VtIur8tFmcdAkZ2d+iSP5mFoxn15cCZgBZ3
SJrwDI44jenowTSNu3rItqBzQkGpRMMzWjSulft/KHVm2Zo3bjT8MdjCGDbQEcWqmGRaWLXLdfIH
oW4TxbPh7Y9slYZwVo9K059Vp5xnMkuPdKxNcih+XlBeohjR93l9prTIvkKc8NtE+CGJVFUxdRQe
96+g5lh01PEkwkgnj1dNtNmBsxhovbcuBJ3qS1BjSIgd/hqVmMouL3M2p0p6969Eh56vS8y81gOA
FEv6wnM375tLA/YquDqcOxV/p0+KxhTNueF5z5cbN1woRmCEsZk3aoPCkMxiED6nIlKazHlO8fo/
7QHdZvyKCfmBuGda5UHwvwYdYNROE2oAovgZfFhYWhQTM4cZfQ91bkAr6APpTZO0dN0Y4hnaZFks
Q26mpDf9qPZfdQzgMkJO//jRhP2lhLKZXFwvETNS05gIxYWXXd5iZfenKEL60JzVrKtW0mI2b8lb
GrnniExy+zOzDNqE98vfXr5tGau4F0mLafy+eJCgOiBpIyGvMLZzNEyI9RE6WDGj5uR1S47nNOQ/
DvI04r21VO8EKnnCYv2bC5VbBB3BcYtOxspENSP3/SazvlXFFaIRtaNxJ8aVXEk97gpCYSAflPMk
pv/uDlIfZ3F/lWrHl0L+aVUU/jskJvWD151kuj2PjyAawIQWZdXp2g+Ci5tf6XrjXFx2mjEN4l+B
OlkJepd8zlWOYDzqYzLosmdtDDUCyvsxlPRP6wBX9PjOEDVsaMs9lvrsTaC8QModFOXzw6HGjScv
XbNLtMqHGAXN2MHhAuBPEeTnXKJtyD+FBVcx2+ndhhuHE0ldIezAOh9yvi5By1D+LNe0ByVZZ9wo
EnBDf7qu3qUWoSNkv7TrkV06cp/Lro4kRCWUdjMViR7ht4kewUyKXvKqcGwzQQYzBhf0KKbonGqx
DGh8tP36QE26qSvLGnpQ449yQE/DMgSbCeoFD2F+WtngJvJTvT7oOv7gotDwHwVsRhIkQD97yCct
0rRSsW16S6tK3p1zt63ikR/nKV8ePYY0JOcsYA6r5dtObyov1xWms+OGUIulGYnEDhtWF2Hqq6iY
Fcx9lOyJ+/V8cKD7QTlub5gyfYanIo0etsb4EnCpasjA4myoYTlIufzkJ5zAhhS06wY+O2drjmiV
6c7SmPpiyPd7X3R0/2/DgcLP5m7xJ/p7S5RGrJvLaMq6gj9uzyr+OfUij/PwCMsGKZiknty3HDOl
M8utxXbfPstXNRAiL31F6vFmMREpKTLV7AZsukSzEKLI0zI14dfsgNgEMxooOwybFqYCX0Z3uycR
eerk21GLU6qo0cjMn2B7f2zwSyxMnQ05KLRUYt4EhddiRmrzqf8O3f0qpVN2d98s4JacJSPYgnkY
a0qRn9X8J3B9Z4MUMLGKBQUJCrIQb4T7RxktHcQuy5CqWEorAHBy+v6FaUPLYA5x26BaHNRMpPOQ
CtMDWKccbrxUoiustyhH4bul1ebZeqeFwqUTHrs2BXR/+eMy9l6xoL2Ue+Fy1/6x7FL96awsLBAH
o6yOX90m62qYbaoDvPjcozfb5teGuIYoqB/dXcMUxN0y48lUHNKJnK4rlSOQ+uEaG4/7hi++uVMi
77HCyHsokA6MMmMs//u71eHiKieXRTLzb37QqjRqo6TStXKAh8MknflfUtMpX3yh9QoNidV57UGu
Q31Zy5I5fHt4/cAB4DpRDQ0OmjHs+P1srQYvhx71U0gis28oYSazk0iWrGNZ8GiCoVe5LdPhE0XU
JH01Z5q+me0/lFj3tJQXgVtFhRU3VDwiVUi/HV7+VtIxW/84siPYGjdrvQlOLX5r8XSZIGpzCWyi
l7HHjt+81PFtXYzzchWnM+7/lhgJvk/sgaWaHL9nE3M9AkHbiMQv0PL5UdI+2aq289djxATM/ij7
Ct+ziZefAujtbXuNGs/72VHN6Fi/Rcbg7Mz8KwTeoBEhshTdniHTiuz/lBvUGz28gYWJ1rQq1u+H
uUJZI5pJkJsCRGr0iUk91D+HWmMFJYNl319Nhs8sXp58V2Cde1LOFOZWTXU7GfNzz1KRb8ZQstIT
OybOa/myWiZ1KUzwPJ7sFMkzBq3VMRr4ByUNKlqi0B4ZcYbHje2/xSAWp3IFqNUNW9s5lr0nLeUo
zI4fOY1T+9A9sd+ia49PhudSGWg+/SDUYdSBgYE8emISyNotrexKime+WbRggz4PmcMHwOfuD484
nRVCBseQmKQ5hmNxtA+q64xuWZMaUiYKX5Q7TY2g0QO1k0sVrtIzTZfc+L6yG9Qt6HM3fKdlTJg3
AZu7VmLjSOGURqMsbnebCIG3lTxFxcMikyMiGb6IdalrRBW/WCwhkKn5FBDGkG2ZyYWSlKs1TVAe
a0rtHndtC8YxRaD7q8cShXwkgdUjossy5hQLD3r4bsatbRVoKfMXF45BGFWJI9QrIASUCyVnNszL
bTEF18xC8ZN2eOemJf4ybmROQo3Ir9Wst14+vX9z9C/ziyR00GBRmY+RRUGIehiOKp9SBEfBLSM/
+iLBwMRWHurane4rTkJSa3A3+pMABNqyF4Ws33Vv+ye59RcO6RhVEteWDM1ETe8PMHsD2iS9bNaX
3rx5thuOo8Cd0XWp1egZRMUZL6pRCc0BdWlc/02g6dfWNiEWjxr1tNp0cALpf7dI80PtMIJTbBvK
unN4FGAsJ8coq0AAp1OQWTEuknieLqQh9X1KNy9Pi6LtBD7iI+S+8MIrbwb4LZstmxZ9GNN5GgPa
Mr7ngyCwwkhttNrouvTBZtklS50Xnfh8H+By0zvKvt51W6cisdz6RjsK44/nlJiQEjMACaIHShK+
pHOluo1UxvCvdRmm9h4u95fwU+zNhiMo6mhMngH7KB3YzeT0LYtY/GZ1uEisgpQIYpog4JIcslJT
IakrfbceuI4Zli5CfXsnJITCRC9t90jPIwPz60QHZQ05lMF4UX/Y1QWjMGOXvufi+rMNLK0/A9ga
I8YksiehSYAMXuObnj9ZNKlzlG0cJKpsYK37XUgTLIU7TGY6jdgcyoFbHJGIqiN9uzEPkLFXLomM
+89emltZKwqeqEqEXgvfo+ru6SrXLcKyDZlpU6+OwmtTh7N3l9db6CycdjOy+ngM6zwZ1Pln7iu2
oEd/naiHbN2/ImG8BJwNwcTx+egAJeCn6LW6mGxSiZs0RCWGJzcS7EzkSfOIbCjz/OCtjt+FmziI
yDTF1kmtaWsJUTO562r3tU8cKAOKqRG1ikoMJEJ//DwOswQ2g4M2XGY7+kQiILaOJaOrULFjM2DM
fCqWx3kfDU3MUeNFUzN5+vVv1DaJoZVv0ynEMALsAPq8UJLP9CpcacxqFOuFiQ56CuKKfydPF41M
4sKWEprhlUhuvDwOnSjMDZKWFDJMcfrj+PwRFpbqt4EOAh5x4QC6OnawDu0ME4wdFmQGkUy7LgHO
oMZDtginJz7pXO174xcistb8wAS7M9+MT4Otle2kyZnZF4RbvtrWqIm06DI5hufwCntPrGEIuuLv
UTjHvEJmME6v3VNo/fCfpdmrZtI1TVPwAAO1whp/jhuKglR9/F2maMgoPgVpAgzqXXMULJQnuLr1
IvbKTgyOe/miJGMHjvCi//PHJbgSZxEuj27Fo6FhcLdsE4y4mZw/f5egcqV0c4Z4xryOWK6/STPG
qqpNg7xxDZ8hSJLPfyZ3milaLeSNt8sbsa6vVzvKz1MBQGHoTXMf0KDFv9WXmtTRrgAXK/JkVD+X
0pDFzGZehtHSGGrlq+KEQ16QeuOHEj/odWSPCRCa1Q+SpQ8zfXd+vRwGSVnNQ5y9F4u2QS92gAjc
no7jQPESNfOulA24uUEmiUg/cDFnuBN5VBpzYUEeSTK8Lz2jEGf0gl5/QUVuiPi+sntLyPygnK8a
jU4vXmrnJmiSWfVQxs5aHur6W9+tVblyngG+9qx5R3J1qUVh3kvrcwN/rNyi+UDTFRkXtj6I7Xku
rgr15U9lgV6VopRZMTbzXb5opZeC9lMu4iGqFe7V2kEMKrL0/L/2PUIIK5kdYpNT6GmIuCnWVVzc
+FJ/BtPfn7kMvu/2AcU9j4CzQ3YeicG4891/53m00K2g4OKLmPTvLC2fE5pjy0kkRP0uWw2tjcJU
94k3nqsEMvgbpZgcn3dq2wS6GF/xRC+BAS0neO/0rl6PDBOdWkEk9sSVMJlXdvZmTKptIZW0WJKJ
+1Z7tWshRrvvMa1hE/hSlqqLSi9nOxtskXhr1/80w8sKR66tpobj3tHL69I2VDZa/Q6G88RBsTgK
fedXVnKAqVs9fw4jhWSmqa37GrGb8Eb5tB8zHeuvu7FDh6r0Q6DI49SN+vxK1Cp6TIrHRocfRuam
XVKx9FVI/nEsDEioZd1t6h3zlYaAGLPjq0Yyc1a6rMSCu7ZswLu5oC9u3cPN9yL4HPBcO6gB+aQ0
2KkMmr2gqQI+CRaSXevDhzjkUjmvkIJJuGG2C2dFSH0ENHi9fn91XJoSxoltawI0hvvd8Socsxfs
vfeXkMGb4yHm7YKSu7wvawJdw5/PeB6Ezo1nZdpZnUy4ogfDXgejYPikjg+QWI2dMdwEmXcLbcwX
o6PdUPIV+aWlVOhe4v9JA6qJ8thBMjfXaDD3DuwaSolam+oA9s46HDJS+4Y/5rUYczN+0hiddmAA
OIkbP36Of7wueFn1ArNVIv0YvGQUf13/hjb4spLEypM4WNZtmU+f/0vnEpLl7+JqeCSJk+LcmEBi
WqQ6iTUZfw0Mhi5bU9O4l/qTuOQjFi2U/jQgvhyKyz5TyxOKbzeoqImwYFVI++mTegCtIXQLmyJz
CNn2UHjI9N12eHSyjLxxURkvZYqqL8kA4pSRTiQNUXQ1Fu32MAeoD+HY8yb0zRukOWPtdq7Wn8lK
FNfaCSdz/N4EC2VUqs/j6Yfrqw+HfTLNgYNE1C41OU7QNM2ZkGt1JAaRcgfIAx9qRCO9K1GpryN+
R0/M4zn3Q2mmTMdAy+UJRo/s8GmfpHQ+bncCvVpT09HKr3pQh/VBbW6ppmcBu7fvcUCoB0iyRnCA
ZIYnxAitOIl2o+J+yqjSvVfbW96zHRsW8bvTY1NBEW6fB2M/pR4da3SSRM96Lz447SZXQnNKn0wc
h88x46TVdExheXH/u8z568DxeVBsYeMNRVR0RzzVnJpBJ08oDz/vCJRG1QN9f5xQsX91sAdnT8gI
2mLFNO3VoyFvwpAZoRpxpBcdO0X9FrV/1pmUbwYEye46rDzvmCn2mBtDQr6eNgmvXPRw/MwXznqO
eFMnPdNq31FNhVP6xNQ55+9Di7oO20WpcqyAAK66wDGuL7UYl9wYdDf8xE0A4XWLqG1taPQQ7xl2
W9F5mLkYaQTrTGrG2GQUc186Cszpc19k2RqO87QQLexA6fWYluy2hvEYbSHm3CRQJu210uvXXdI5
PcLm38yoCn9Kf7k79Ev4wE88FVHINEWiF/RU1Tpz2+loLNK9zLur85c+1SluLM6bpAn1gF4bMQbg
G14qompkZJcgn7HfpnKTtttrAfn/wwHWPlKSJowoDEdQneZaeZPmbfhIMDKtahrA3YbVB9Rk3hzC
SoqxZDxFQc+GNhWCCRmHkWoy+nFHd1zWsoiBXzKipOhDml4b2gqzO5xMBBhbz803nP4HXY/zfW0p
bpChVOid/nhq9CgH9qXhb5lrQxIoRXH3eOUOtzUYZI1xmgdObREEe5BzhnQx1kBiziTjsncA6l5j
/E+tPk8d8HTiS/3j6oXwf2/s6Nw8mq0zVoShHLLEW355EB8NQyrgIMoRnKM1odiMpXrjFw+drTZU
PbguLaFsRuwX6hTPf7bnF9qJHS+GMETw2Xnc5xGax43tYXmClkxJgbJLyU0QnGPY+ppl4wnNlMCl
LxCtgl0k4Xu17VDv/2H6d31mU7YDOQFFG/0xFGma+qsrQcQV53I70udMMo+nF44EBoqvAfWhKk9x
hUms6HIANt5R5prdE6roqOhopTV/IctqSL+kMtpJx0d/7Ccsy0MigyUDVNHohrXRiDUcdTGsbsDl
Yd/PGaUDG2m0wKQuJDtavp30ltHMNBDrNvi+rlfZZNnE3qnhfWLZD1Y+IE0hDFfGtV6GjQBtVCil
kktegcCpXQjt0TLX9FFeAYXb3LI9CtzN3n3gTFT57+Owcph6wx++pXpY925htNjzo62eMb9YxTQy
xG34pMP8V2tHqXQwdvKyzlE+ocEjrZx7loyvn2Q3rmBb5jHARXfHcfcObetUkk3e7T1EuM5E03Wr
ilCcwsuSIjzU1CB1/Af8YoAwSz/tdt0wJMgXrDuDYaU8r1O99RRXnZvg/KjDCffTXCf42pMDzdmB
yKsRYQlxEXdJFPovlyh9umlJA1arP6+s8GhHBiQUdQhEyYpRdmReVrc6au+lPN98MJAdErdk45Pj
seakriZyxzsjRo8han3kvZGmQaHYiX1tubYXrQSS50PJ/4pAR1POS8K+kowpm2DxjH4qBTKSowLE
vLUH2xxKpvF++jrUMiZWqTSZvM4ivYQpx7r1fl/zykVkhpxIHnsl3oqB1Z51Dr/scyDX/dp+/W36
dIy8ds2bFmg1wCyxyc92iqT7FQR5JMzhzZbPvdJkedPwwP0bWG7XK2Y6deXW1pKFx0cr4zCwQ3EE
oiqlwsDEomJ3s4OJB0bZEOU/AMT/VWLiH6TE+cOTFa644564q2AjC93+bKlxzMiAECONEmALqb+D
hffVKtevajoC8UsJelDkJgv2eM3Rhv0/Y10r67sO8DY4WkUFOgjwwFQh0zjmIwKQs2FJtycwmUEy
FJ1tU0m5x8Eay5qsiq5v33bga3NEPMwLt5GS/C53ZWXvxUF9ZM2hAfj7xc5QtoZacnPgH7a6/CS2
NzmmCFLquO9MOad+G+ePysZc5I+lPdecLp0+t3QX/XW9m9/YBPHpw9iwW1qzUJVP29ggSqUdPpcf
zSPcZO1pRvzmKWstwz4OpGWUEifbL9dQCO0zdbbXHkC0pRuhJKLQppkszf3D2pIhvGXGQP2J3zds
vg4uGkj0eO+PqqPINhxqSRcaCE+mYYAZA4ROjrraBqqfRppi3UwIUX4RH3GkgOWnZl/mBpLGtecO
jy4+0HrKPUXAfDfYYTIf+j3jzoV05QYaQcNz8pALh/RVXYQmcG2Mlex3+LLII5rg96fRMR3R6QiR
/ieAa0NqN8iDkPRVSMStnkvoDIxuDZxBWh4z92a5CI9EO5RLoHFGxFk8B0lgvrsCX079DdiWIPfn
4MGH3p1WwQbWtRQ4UT9YCWy7ED/DGaQYb3plW2Nv+lciG4vdtYXY775ILQWRCAurqOR0UBBHU1aG
ma966IFkhCL57yqAnD6n7B/hYwr0gJhEJO24JKnkH01Ns2bW/7CQDrUC8Jx5mql9rSKo3QHFzZLZ
It0pQNQg2zWj3FV7E9Tr4D5CNHG16b1kL8V1wJUqXotZVUdOfOJ+l2IQabEXhNeoSeyPIvkVHkNv
rVSWipfksNcRiwpqw/PWUxEJxh/chAUbVBXeXSiiAHWf6Vd2aWNPEzthJ6m7nH5IeuQ0Lnz81tCv
4SKUJ7un+d2wYbBQqak31tPdWX6ao2vNQoQdDshWLQaYSChYWAcxVHhlIgIl7qo9kqWbu4YWTxW0
ndN/GYLhBpYZ59TeWC+y4Ml2dq7lzJnXMcLl+bNaiFX3t7Tly3ppZtlsDc2KkU0zWlLJ4GZe9iFX
I2ykixkYm7KT18U7mUvngyd1NrP8fYuhmce0EPLtX8aPGvsxKaV5NfN/e4MbcCmI5bGMLllN70ND
NG4cKjbV7lE6BaaBtwpGl7MmIe504h0jhdAqjXdAgLeb25StRKWRfh5aiiftVZPfdxgJS3a4KxPu
ZrzUG7nwtwYN6jmgUWZZ5+GfrsGFc6Uh7t8tcadllM+s/sCmJCNknVvSAznvlXZQIAAtDDuNBf2m
q73EXItNfyg4yWIktBKGfMMQeOIYeIsk3ONUSPvzo2KYAJi7ef/ek82SbRn6mNQTrEr5RZHFQc18
yinfY5CYeNpVfcATZzaUvXC8xpayxv+7LbwQQieDt5T1+svvrMEMsqBiVI8ROO22iyCUtSXl4UeW
vG6YKLA/xSP1f6dnliY4zUoqFAX09SyIUckZgf+0bNycJi+Brms/9xe/sux4LG+GPbMXDKGEh/I7
2lKhApneUldX8Ym9Yh3gYtlUCLHpDY5jV9Iwfn057oHE/BSSJKPGUe+k8xfQB9y0QJkdSvaumIPS
AbeUnBfUJxqHXmAyr9vaFARLzmiejs1NvtwCHSWp767McpDNcC2TjPG4in244313cbVdB6jpSAuP
xAw8elaDum8XrWEJv3zDUrpgNch52kXvrF9184SAW55EHE1zsMYL2tLqwuHY9k4QYDPG63wmlZEf
5Z3lo4Mw4rwEvQeOBvzo0t5ajrCzlJUQK6+yZX1Guftuym72ki0nj1INQHpIcmlTt/0Iv2Pj8/fU
6PaW5PqGT9s11AkKenNUrpL3dpg0pBo1s0ZR6G7QHU2A03JOX69/zp1X/8mUCLl8cWkswf7tzh13
U7/NnGxmQv/fVHaBR7YQGe8aDpu5UMS3JNohucYjvB2QgH4eDPOZbXUmV8EpuMDyGxH7NzefN8c6
zUL4GhHnXYinBU3g7R2ZdRgXq5t/q8dyTkqyS2jvyugsTd/VcZkefb9EU6srqvSY9LFwBVkGcV26
SL/pVEq48pWZ2P4qvcZ0+AFyUSKSYVCNUVB7HzxwEBP1baN/xdouWbr3+Tg4P51Y2Id6p8D3n7+P
muPfBRoJVs4lXk9xo5rorkHMyTK0lmraZxAHlH0QsAmA5+2zT4xiLxrfurOD9v0HSECXNHO0YCFC
OltB8O6QM8M/xW196voxXbhujq3M4BWb7zKZaQ8sYyacaJyCHmwQIqg8J6L9xiUldabfjD/BGQYi
opSMkUv06t5lTytoejxnZerkSWSYV/1EtEgFov6xI3jW53g0Zlr71sJwaypIsrNwesPKq3wI3Y+L
QETbui7RTM16J7UZnDioAxSxZCYpuftxFnMA5ieq2Gs4SNTSGCzXw3sP6hizkDGOZRcEYtYEan5L
oH8o+7TyiAKycrVmQlrf4aOgE7yv+0pEvf9KYRSRr4EqQOy0MSr1PT1IvIcMfdjSKO/mgXQ4rwnw
B65a4nFULZRcZTdTelS+Thrbc4qUA87VdWFGQz32bUj9tTb2m9NNw5VgaPDwKuEQpxNZHFs4H56M
nLkIz4II+MmulhepUc1+wxDEiSBXI7IEU/y/6j8eWNEQH+3iaA7cXvHx2iZHJjogBMc7AOObHZoO
z+ZfC/Wb4c2uJ8biPMyPV6DKyyK5gI/9MEp9Y4fA3BqIXDr9ik6u2UCNev5sRkKqvhrL3T75UDLx
2a1z9AFsio8a4Sw8RozQB58ilRmhuLHkKFIW0ZNUuQb8rrCqKbZa9SF08wGhRuG7HWDwUwNl6yaN
PdYv+nk+gJP7YoHeEZIF5CIKKiZInphjUQXK8QefvZjggERveAoWutWEw+h8mlAMVkrHoxd/DWfM
gFy6q7YaQDNPj9c2kIh0Z7dflGHF+Gu5I0oQS1bHD+USnaXp8Cg4gKulhS5Fz7mzJNgTR4EtJkpv
xALsEqoJ/GtxlADzSYUhFRsDmRgRWVHtsGDI9422p5WNLIgK45+pLItC318y8Q/Fwlrp7qfs05Lu
iUBUkvihV6r/+KffAYKP08s7nBq4FAG4lPFmicNGc5gPWcMAqYwtqMoKtXnOMIWNd7G4VGlhvUmq
zsJdW/zI9njkVHaj75X9zF2XZlzp5n2CG8mMhqu9UbROf2oZ+k6X3RRTnbm3QBQPxj1NgdaimRJN
g88U8eAlAmDXeazBQ7E4QmrYyVRU9AEiT3Q0i62fXNgcpet5Umvg46GyKlfAHKvWYIvAnwjyyFwj
SKP1tkPboglTuN3oS6G7KQ+R/BuVkih16v16fMi5h15H/65w4RKa4qAnbkzZanG3tUsKoWV0sdai
RsvWzeJiaYCtCCR61zMx2ljfouKXhE3hPNXQXt9fFkp+aBjFxKB2YDpk0LUtRdGCVWPSAvTOdByo
ljBq+flNuBwzllrsnuJZDZNyj8ilAF0+PkIfXW4RTfMses0z5qix1Th5HyAt6ABo+5Ov+1GBWtQ0
V4hJBBWZGc99y+CEu5tBdecFW5ulWhh9+M0nZYzdOunXiKdVaYoZTAYC6fSUB1edtrtnnowHHRki
lLv1lMDeIZWU9clXAGc1cebK/JTci5wVJBCmnLeZTaSeR2dok4ahB2Rrd27Fm34gY3nqZQNzEmft
fUVQIhJJU04DFY6ny2hEYImq3wS3puVrwD5fEzaabzIP/dkXkKHnGoe61MVBJqpEtziY2xqoOL4m
Xr+HxaIrF9WsLI7oed5KP0jsHN131RNTk3xPy4W3pAbZv9dhALK5uHSVqL1RjYMYHSySBR+MsB34
tZl737c9QyQbD/SUHMCO3KLicDRKog31aa0DDdqtrqBXM7Kjhwu80Qa6dOfErO0OnKwInpBzBYIa
sWX2yrXwPYFgQbtaJK28LqfbXNQABLfWniei5bb2GA8DmJpZMA2AoBYO0xKGmpcCBUWwcPdoHsBo
DGwQFlOMLkewVl7ZmgpHp/ZMoqAy9Rk/cjIPH47dmgbRc9xXso8a5hiRO70oI8JvvKqrDodGRGH5
w/kVCKXXv8Ti09A2RFQzKQ1ee1PYrw8dvwD3iZDX9BK8cuEwb8qoJL1w2WXdjTJBIvunOHSeQI1T
2Vy0a8t2QSZtxfV/UlKbotNXHJAoSFu5/Kl6WQ4L592qKhMr2ocX6tvvAaTRjBLernpNVx0CsmXb
tXcG6x8yDMhuYlZboG/5jmt4fUEkRvopvP9tYu7cxAeGi3w2i7Rljen+OHB9h4DYtSwKjKdRkvHX
H+DUNGxo2AAhlTamw0N0mTY5uICJ84PHbCD1NPzu6kU4Ecr1ndEfNCerJhJ7/25bwK3fgu5n0tq/
NKYjAOBh0B4FHf0ODyMlWlump+XLnmABVncoJKN3OXVjofYjJjubEH26MSJyFn3H3s6vYanDkhTG
wpqM4m0+r5BFwnk8bT6g2JGObKkPvJ6Iyf6djo6vYZzJ6gJ/3j9AViUyfvlGflhcMKaZwrOmmeZ6
Qi00tapIQ8JmREDCryi2hgKQhGM8ZcLlxI65RZ4Tosgw8v5RALtK7R33Z+6LzPGAM5ukSNAqxVNV
IAid94dGbLbtmuVeDFkh4xrHozKUeNP2XL5iabnYHXAAc51McyIEunn4u1tEOv6z4xjT0yMm4LUS
3DYepEtU2yxF0fTnbEj3zCWY+ZK2e2u+CahO89dUGMOdHunk9zFjTVc1p7DqBaI8kAUlrCa2UM2Y
6PzouCtn8tQFZpoAFJTKTPhmZpNhwLwSM3HACZZ9iSmCR+H/116JSrC7kzhO1xh3WYMFTxujVeSD
WADY+5H3K/7kwkAo07RDnchYtDC7mXmXDAbupzGOgQ+gP7iiAamrALTWvjDE64D7ZHHKfEY9qB4e
qNCQwfKU83AgENqLZP9RsIQnC3xajCeVXql5ZEVty6l0Os1E5Yyhy/cRlt+aEoYF3TwD+mjlSFoR
akRWY3WZ2YMteuiZGJN9dGlJk1DZneYIL9BafSMqjefJDj1xaxITe/kAOYbu6Knm2hlf2r4KPzva
nDcMWlSmldg70/Zr40jL8JxII31O3LWRt1BIWczHLH2cccsvjG6NOBJi1fwyDuA3ybWP9a8QK93L
Ls1JwQX+IG2bHHy13IQmEZOd0ZVjn18VursJRAMtPpoXw8N4DqrIIB/FpZDFTwb8OfJjwiADj9mC
mRAthAvM2GN/ZwnpxQS0Nnf5HPhbLXuZQXVwtqPA+mPPJL+osjVnxj6sLghJCpVvzPDXbjwYqE8i
eWBlLgBATOVWPhe4v3QvGiHvLD2n2pQl9tYHGPGNpNrmrLfjZwkJRhMdKkeWxwYe629TJW5tS/5o
9T4hMyxDVeZbOSjWVQG2CcG9PHs+blLTFfshAmQLjCNS0npSzI83nTWum+CCn8h9NRh0mv/9kJ1X
L/uX1Q6egL+CkhneC5zN9nUV/ph4G/nYBSsVtXrzlGxjzYNjJXnfAdfXQkDRpxCBeCXMoGyXRrxR
mGrOXUzOdKfgHz+syTkaobwi1Ra4UrAxl2j0qis4HB0dRiPfAwYhBePi8TTQkoOAEanlS/tEcUQx
ovpvd13w7O0c2g+qwgB/BW7WumNPDego8fORUaDWQbnsTL/iNbuhqkhvdK1kEE3e1IeOftILFVJh
HKPMyJItbtzglXz3zyqYm9B+lfyNQsT2OeAHPXAXdkCl160e1uf/Q7ETLqj3BfbRrJFkmwqOw/Ye
OPQtnamWwg0MBftQSXOj7R+RCovbGfQOkUclnNjZS+PFwxok+XUBa2PcaxKDz4XxFgAs+E6iNLk0
CZMnO5udj0O0j7mFVefrWbxIg5RBXWCty2DAH+MxUGD3GycrwXtDJpG9kN2uu0dzViVfoSMe+fUX
+veSGFUNOo5z9HiGsjDNmdOEZfl1B2PLGlNjxtnMpHqWoEjOdIIYvUxABXVSJhAtqdFdZxN+MlDB
ZZ/k/ENudw+cq4hEMeHx4Lnpvl5aADEl1K8Fac0BSR+zR22XuNAzivMkUXqh8gKP49Xd99aOQ+uI
pXw9IYEpJJUMbQttqezhTtB3ZW35oOG4WUrD+5hHixg/nh9QeBvjDgiIZN/gTb+h3ye+ab4nHrMD
FI6Lj3hgFPArUlD7OOnj/plv3pjsXHepjPqt0SOdo8jW2aUJUra3GGYMFDqstDAqJCXulTul3fJL
BEg/gqUIVkz8ko/ec1iGj/AYtK8A/UtISSRIgN/ZuJx+3UXk6M5d2gX1I5/CtT0a+n1SGRGio5t+
wdU14cyFi14D8IPl3GSsf/4jEGoRMqbDzVCSH1J9JnxtyQbDbUU8ffVFfsWuKnO4talXwg8GmqUY
/t28AOCnz81t/+fFIYa9M8Bm3imQvuUSbQvaHFwqFM3iDayNFcw1Xrc8jBhhaQkQcvL4ArTNmflE
mvszEycnAhLxhe3oS1sLdvuA4Gmlq64n2qOV5653Nvicv7Rgxtg75nuTwL30g/0LfWS9LB1gDZGf
MMC0qoZlICIvYqGs7sNFUIccY3dx0v2nVLVppyYEj1qgGipddwJfNwwzTwjiOm/0vgY3ayzA+yvh
GsnFKxJgV9Yx4BRv4IVXAyNe9lebue39Xg3m4Zpe5wBxn5LcuTY8ZWkJfPQeO7Lzrs8ylyXVu+61
WV2/i1OrHOkrVrZOVPpayaBDKU+xBYd5b0fZZKRGBVtTE3t+mzqBV5jS/rtMdDFkBlcwnXrpEKIJ
yc/1jyVIlmD9W7scNxJZI0ZeOnb38fFOXazbb/C4sRaHDJwjUJc5qUqZB5q687JAcM7UnlTiFvZ2
R5aaYmApb2CuVj/7Gyfu/2lOHh8U7uLtgZD7gE/dLr6LRJlSEDWfIi8tnI++bjeCk1ReRJjHGY60
IaNNkYhJP17WibM+LyACWh7212Ds/jL2FF31i5THh31oHhP5gkEldfKUa7Z+UhEiC6cK662br1V8
V96w+4IYFoY+jmCNFoF5kY5yz16ppm3zJTCD9VI7d+g1RcFBc7BvqhHe8XzaZaojItNHkpmRaPLZ
JBuXOOMDK6oa/vKQ87oZL7pCwm7ZEKwAfJ+JQmH4W3Ik16VW3jdZ1UcwPjeXyB3XA4heosMmd/Gd
kq629/PIXd8ljWrD7PmZh5Fm8uguGJpIdOvKJZAMWfNXLRQDBmpNpeblB27sMPNMCSTbImUqnbAi
VNxbJHEoI74CWYhJZYNBFZbl//bVbS/bjdJnAo2nJnk0X6EK8IZPy0r5KJCSZhbTP/a7v6W02+IY
A3ryGvbChkmXP3kIIuzdsSZqBWdY51IqYJU/ebHcGWfIeLt3KlC3S9VKbF8oyibCTfOlLHev4YRV
LUZ1D/JwW+ppi1GPAdUb7wjy1XOZDVSakijVDifWMfFdeA7dUwky2ELfDNR25hZ3S68MZDFyb22E
brPJGzpV4hXzt3rhTcx7ZataFQRivGVrgsarsL/Kj3/gtbChONJAiLFjHrMMNxP97ET3QYZftPva
su+2OAU3WvVUCTEcxmq7H5c0bUgp4q7zzrSaOqHaZcOzsvjdYVt/TxCDzjd7U2x8Tg5mm7Vaj1wq
4AZqmAry3fgNCJchJfMpAezYwCTaUnTXUEeU7Q6edWkEFQVqSFFDaSk4zkWqtMXdMifYb+9X5hee
jzDejmB8wUZSNY96/1sdNV6vTTJkLMQqeEkpC1+rBu7QnH5c+qIv2RVrko4QUqzh6HKkYvrBojJh
09Z0I7poxvZ7/omaM/aPQ+oUMM1XybpjmO2zDIlXPUOQ4xERpfi+xQPX3qS6wUnc00QNtx8iYDCx
0bgHVY1Y8otWCTwv0NSJDPZzAwd17zcWiQdEyMG80rJG2K4/I5J9fpbsCXDxv2Mgil5DSUaLoa/3
muDAj9hA/tfZ8G3XQhxYM18kHRWgsIcXNUI9S3HZC9K/Trt1v/vv3Lle0ZIm7vvwXQJUJZQGS3RV
rDu7rmBeHTiR4j94N+KrnqPmZMWtRzRHT7xvCMJd/+SkWEQ83WoBstZ9exRqxKotEU0pon1dO1B9
G3fYwZ1mXBftC0QPKAsYECctaw++jfZTkp7BbbwFmRrsJ+sjiSqksWXx9uxq3VwJefy1+k1yxkjI
/Sd1UJuOQ53ho8d81Vc3GgblRHhyaW9rNsTCAv5ReXMUMRnrN6egUvrFfnA9QjB6gehXOJxq+Rjy
2TICt3E/0hzIWpIn2XXvPrJvbdyF5uW0w2XxrlKhk480B7sDhMfQav6zVlXj6FmepYxnhNIS0r4c
tq/4ZMRY2ke1R92msPM9luJKDnY5gYzfGtQmzVN+JcWdYHmFNRGPQJ3usG45B8m8D+xHDfjILbfx
nGhtO+6xMkI8GX2qQTH9t55Y1D93BfGuC6CQIEKquY7j+A6USlQFlpyDlz1D8gMf+pheZ0kF+zBU
qbIyCSDT+vuf0QUg55ApServdrQVxZqvfSMVDC1oPiyf/mh/bxcUz05td1zEPm+Yvz3swvC8aJWL
YBpjZnCz8qKsjEa59zPNJOgRTEeNChH9SFcHjDf4QIcWfJ1EUoLCZDnw5C4Dm7uLnJoSP2yFsGUK
cbpKjOYJ+fcxn9mHpRwihORSvugJt0ZbGWY6s+77GJ24gPpoO6x6ACjmnSExC5G8uinG0D8yMcGl
AhM9nQuXHFkyj+34JsciYCTQJCVPnzauO+jE4F8lJO9LR5Cs4/ZLidHVAU/pnPWAoDRFKxGFCWLe
FldG+kXyVbLtaRTvd0EgkibcpA1OttqJvkYPp82MLgwgUaV3ylbktoVe3XgK9kKteFagPcCjkFpK
x48YP7Xx1LaPKeDnGB/BszjefuC3dqNNoD7xhs9HvNXtppm4xiGl/CezLPwnB/PJokWkppchnb/H
k0zfIYk9yfGwS7TuV7vv3QexorFMCJ4rlWIT4IqOImnynjvyyG5ba70GCv4BoLR3eJlD6AbcQTqM
/Yjw0OSFCM8OvwEG8Ug2NrcIKgmPhrLKFH2Qrp54bFJnjS+um9zbF00tVksoJOO2tcsh+wCdQXV+
fKnqKKKJQ5jfbP7Jbvfi9mAnrXd4gOLAaSqciupRH8b6CHfFZ2kNxdqNc3EpFCSoR1prodAyBF9T
hNPeP11kcIoPV6yHyiypJDxL793VGPtWQwjAm8BVM2L7b0KKYE1LPsDj/HtFnjCVWQPfAr4VoOQi
qFC3kUuJv+31PFtwQHmXh6srqixxkXpKfBitpZef0DwFYKj3GlOnJwRJUXni2UmDMTgjvTQ4nep5
91aPkM/vZYTIcPvfm0vByt/zYnLGfiUYxZ/N0HluDdTS4+WfzEu/Njgjs9MyifJXJeDswq0EQkrv
rcyz/y4goKLh+KlDYDhnBV4YPVpuUNJuD3EzCaj2qCSgjY1u762vNJGIjZ71tuPzIoYO0KqBipJa
wle0okFuZhtOcHqIkhII11WqImoo74cozmc3ZhJOe6koRS01vBynWOOXj4ZZumtLZ/0J/KGkFOiV
HftTVy3oVE0NmBmze2rh6UTqzesPIc+ZgpWcD+070tey1Lc2AC+wctMQg3yeWARePEZh1SNYusMy
OwKA5DNvpKMKFaItyT9I8cMHxCrFKbsGMmlIwSDn3yO0daXamaUce8ww3TFpKKe9Vg2akL1cvy82
Vlby31bHSenLwY/W48WRnmY+7SugjHirycEOBQG+ELSbF5iwGIZjN2uuaPN/J9kjOYg/b1TVU9JE
yRo6d/aM7U/gh//bFJz360G121wf5Q8b8GOsw1ECKDCEVcX5dCPOZHNgbH0nDI1vq0/FMX9EtCF3
yAoKe/j6Eh40PVaopsa1e66QT8nGGXqMjuw/wUNgQCiEL84/XJxrpDuW3K4sJZzN2ax1BjCcFOna
JEQoBC5jU/lgWKcMIJ1Qpk8ZyQpe0Wu1s6+2zyqNevDBhDIxMCwmIBeRzwILpVFXdhAYZ9mnpT5J
B+JJoA3BSLzsa6FPEoUUsgPhqa5hcVzrE002CFxMXzA/egZ7eyYC2br6g5DjLdgiedqSXrkwrqIM
qXKYcphlSw4twTjSlI5/kID9ww5k18Ugq7aRd8nO7x3rvd3BNkRZEEgvUgh7MqkPudi0t0WVv8fw
HIKpKuKTmQ4J7jr/QjxbM6zK6XcBn1YDPAo+UFBCm1WgLBKKZk2dUlz9U+1+cAUAdtfydfbohxgu
hWEcNZ/7B0pOdT4OglwlG1fLV0fH3rSSJmPsxRdOlrpSs/18xvT6xoI2TB/r0YqsHwHtlaMc6NSt
jwO19d8aHAGqiZbJ4fcw1KRi73JUumf0ZXYO3y1fBwRT7tq6LPNw/eNTY6RIu6CI4VsZ0Hkjev94
1BqzDzvXVexByARuHeWoBlbl4ENXC0tAP5Y9qixZ4+4dbLd+3WVawxWdOlOXY+9AYx3li7if7Ow4
ejlMP+NUL09VSfJTlBlHFfjzDy6f54AeBWBQDguNNoAEZg+f659H8+mzKN3UWbxgOpGK8n6M67ef
Xsw4WXFQvYpMdyezkKgvP2EjYAKPOwEbQgTGJuRzEwYpyceub9iPMf4IdqJnRMS0AoUCYozXd6+x
WL2ixORkSCdPhzAsz1O7+unzznMb0ds0ctePBUrFj9NOfyq1zrGAQCPdtStruvFZ7pT6A1nB2IDV
yuhHo911EO/l4Rx6st0IvywnCmDZP4vkdXsvmjnftP3+doRcWX7BbO8D9Hq5UoMrFnA5I/t/jty2
gaXc6mrUoTb20kuBLbTjdtHnVA1VqdeHTdjC8+2QVcMtwii7qV2YQseyy2mFyKWSfV70BrgdO6mH
d2gL6Ox2tLe4FFZp7SWTN7f/u/Phc3a88fBswwP2nFqZCoAy8ic4V8+kQ2+HiBJCTgKNCrUoJZf2
sUYeFk2mwdqC+pF/suwHkkSvzNE5YIYwv1gGB7LECQenxJioB6DMRc9u/G2Aswt2ItXf0Uq76/p+
XCegI2kYpDRdz+EjaXNu5KSH6P/wmn8vWTfm8Kka9LxCG2w4L+9XGDkd4xBrirKbJfOS6Lfr+q6p
iASKW+LZZ2V/U36Zbc90NWvoFCa9g0erc0Yyl6c2W3g/c4zN/0vjWKHzw+c7mRMF2f7+jGPz1cS3
ZJtGwlf9wW4JY8Cto7NwV5TKI95wwzvltwIV3ATIR+NXKbWsFyrTBBpbLybjUEUQ4Z2SUKjdXKiM
/U3OVJ4FXkjb8hD2sHvU5qst3DldMp9n60m3lPI2Y3r8VxESKwr+Ne6tCSWcB4mPJjrvULqxKB+U
Lovp6+etpQL0Cd1sl/uws8vIsh24uXrTrrN7zPFu7rDaAV1Dwcxo/ky9pe5uO3DjGc2kbFd+67Kb
Y1qYFt27XKCtZdr7qwqJhSX6G/YZoOlgCRf5lvhe5n2v7BH8n/kNl4kszhsmzsVg3kkza72Y+FyM
L6yVBVAAlzpEnFA4w0UED8wvH42uaJOG48L2/8UkTO7bZzcObdUkxCKETjkoDNTRZ83DvRQryBZS
vjGJbtfVJXKwTD0MiAU2HA4okKs1Gj0ZSkr+ZZDeJkhmujhvsTlGEaOwo3JuevNsSYW+MHNYT5kC
qbLdnvtta9S9YzEJRQlLHzFdlkK6McXdFO+PKVjurOzoqs4tKbQdWZdk0ZbS8Tt2dxIBsW0EHa3/
hTZuidy6jrci7XAL3CA8JKa1OxxyvsXAjBfNzquSxdGc3IcbAWoKsUbKFGlqNbPQo6PHajRDYYxD
d0j+7sUnZteHZJxaWj3+y5uzUS4sa1iccNrQSpoAwW5SI6GA3QyMr9zTScKU7SksAsoM9gUkk2eH
oZ8LCrj6iVYSDBisgPUCKqJgU7FLr/ljUW6fwPi1hQJlA8kd0R/uLAC+Ny2hIxV0DdWo41A4esuh
nfBmdJIpytxxFAUaksBMsS097vSgN/1PM5c2Bv/Ww+k8Xg68TcuYPZbOgPcjd4pKtxGGcX0FMFqU
6skXzflsr+e5IwefSLLn4COGk/Icirr1msp1wIbuuoRjc2+/3d1WWdHclfkSLyqbvngWHuwx9THv
4onD4PRMqEoJcfY9jUpuErjaZgCSHtf8BjMKzIZELaMGAJ6gNEets4xLuKWCdrDgA2+a0xh+ihmy
2HHTAX0jZAxsZqs6QTRbZldHG5vkdW5eA++wxMrbqcppNPBAhP7qbp31ndspRZEYVu38PClcLcty
6om6Z5Q3e4EQdLT0ZX6TLJuzYdqPBcI6HCaLpdo78hVZiSSV3P4kw7bo23wtTEN9IpJy+Ocn76Ed
cipe22uMWcQUljUsUkB7YZYQ+zU816yXs/N0LqvaXXBhPOa09aDFe5A/awOhujpkX9Zgv05apHzD
Ft3U+vNyCMlrSs7tH9BrklYUIaAO88b6yAHnPYOudBmIThSFM/Fp6of9YK6igXQ2RnEgWKPXIsPp
IyDG7tDe9r0JBLCcughfwdX10O+tiWH4ZZU2F67Qw3oSN+T2aNYfked//xKhkw29TeTY7PIkm65X
4vEoaG4q35H3UZ/27yLlKhy4hJ89kz2hkOdrbGdVgrhvMtuVn/YUFffW4HpuQOEosO6fhd3qYtOS
2tOTmM3nBCicSirolLHow0T3E2c179IWjlzFL89Y/+CaPhTUUhmT930dPTMHwOtEZHPyyIx87ZZf
8PNLmo2TAti22ALbhfGTtThS6nHc/tF2ea0YbYFveu8VvwJDehizEaTdZ+P1UqO+l+7lzw6kggfM
a/ijsj6xPxx4m1oj3mFJMkUGC6l0GxEHuFfW3PATRsOXnHDvgh7qQMp/odaQuUHdLtpEKSngtxVH
QzKh6mqNl8i+1D/CMojmWePx90uQoh7vcQdcXfUZdsPs2bHRtptKqAs+rRk+xtRZqVRPJWQlxewA
qLW8SHv7YRtRauMSfhntlF58O5PE7YfZHuKSg8d/51OI7OUCgDp6Pe/VcPZ6fchs+mjUkyZmI+Rl
1IJ5PO5sH6UP3W9iRNmC14Sgpz/DCH+TUZK7GkHo2uZt1x7zZHCDt3u1OvgIQ5fCSlYw3n9QIfXG
d5qVb44ecsRVpfWo2t+yuuREZOgnFmQUEXNMFCJe9iyAiojJuuU3E2BCfxVO84Sh9ZvRJ4xVKUx2
ms0EmlNw2372bacG3hOnOQuNzkjyrAPZsJZC2KBC/U4seiQK7gu7o97i4IY/aigeWHrrCmrOfsjk
LCLsFdk0myvlbkOlnxWk5bBUXKqr6YfYfBUVH6jtjyZtUSs3VLWvFZcynr2nCzzgFroK0tH7vQCX
7r/m78Oe3RRPJn6pl/fx/fA0sEJBsCdO3HQW26jX7AA6rlVOZoZ+mfDasARFfrYneERQdXhf28wX
upsGLdh9GtarLy8K2ims7xMsakeICJK8YBKRbPT7rdSp55qCGYtnEdIYLEfeQ29CAgFQK5ipHBzu
FgAseRkLvdTI9XosrAlLtkckGKnvPizxxhN7mkxAaGNW2SOIi8RGarwBlCE91xhRg/2t8IGQIDRR
rYxN4H4bSHz5XnEnxfODAETlgnRpw3c59Td+/qxWN9OAiQGk69TDz3bC5GCoGJtNFINZmScF37zW
RRMTgvYCiNpjuojzbIwxL+kmxt+8DbRn3sW/GD4Cj3aFF3Iqk+UtPm36H1/+hWy9M2RaP7ZewsaN
bE77aMFwKIXkMoUWbGYO7YZnniBW3y8vjUJ+3ucc5T66g7t45omdu0k+R+dueq/6CGqH7LMRI6WK
M+Ni3d1LgykSgqmKuXofWRLqW8DGcMwSxQs3rVZb8Bv52T8sEO9qEuupCcsNdGBeJP1LSawMHMhG
ugNdBr+edgpXrJuE7VyTNowixRz1nDqcdLd+fBpBvfr1FDovXkXyuTsYV2wMowECPTL4u4OWtF28
D9YRJ0lUKjVnRX0qwnroueWmscInmHnLKFf4Oo16U3c3tMgeffNePV2ya+Q/oZ7p96ulRrzFw5o1
HhAEyxuge0f5XDka2OvGipp33nVSHoKRi5nBPOAEJwtOWZyxVouy/m8yB7IqCG6TwpU1RJbVV4A3
Qt4PCLdYqKivoWnmF+XQdGUHpiGSlv66sDSVjXOVE16DZHKxWTrzhBd6N+z1Xq6zFVLmCC3LPxkN
yM2vZ9ah7937xug+UQ4kYE1yLn3k9O0xEgEV4z/8nixdj/snfVnLdSEwqq8xRnGYhlAB0MsTbueI
Z15mXoF9lIqD8IHlWhohjn3fW0k7VXQlw4cBf98wIrSdxtTWRLc83qLOXxdKm5/Gj1uL1hfN8z0y
8BANav8b1qX1hBG5hSEMBszQqQJaTHWZOLizQXM4Zln3/HyAzlUT7WVlJwtqmrJELw6t8jpzg9OH
cWwJluQ4CRWlL0IDUTmfVi0bSR/R8bs2dd2vinUQsb5DFUZU5xkkh9VQazEk0/oDgt8tSSdveg3k
rUHRjBhwlGB51hqxEySNL6IUTcPzAFSTrjn6fj/xs4ei58oaOhbcd/AfCxVSNIXp1Zu+mksAdoVE
Za5v4P4EGl4OH2zNL40eKCHXUICBhe7jejL+E33M9TZcDc27XWQ4zXqaI6lbtDbIGBSIValkkgcy
Zw/3y3KMFCnJPbWLab86ajY0asvZogShjdG+dna48SpU79M7HyRCBp+WIiIRLl1Vbwz75BaNkJFy
2JA0lTzERb1RTWdYKwoWIknllUJAVuY4+gcDhGFC6pAvjjquVeK55IBBm3mJXWTt6/lXVGQGSSv1
5uoTe5GPf8K8iOmN+nf8hSTKIFqCKoG5apOOIrQ1SIhn+LJ3HDaZu4POzaddu5v4KgNHWhAfs6aS
+Vdw77UiEGbd13IZuTqdiNKHzhfUWQw/4yRTqRnRnb7oEIiAJGlZcCUn3GZWb69TmXraBzq16Eta
1Iy+Tomq/Mnd2xJYl/R4qVWw6M0X3JluqcFInp76K01/A2g3xFtBxQ9gUG8dlCZGCxzTdqoTprPF
pHorc0tEHiCWYgnonS0YG6S4OFLNqkpVGC2heSey2vO/AhFWrdbpUKkMZDSJ98HFwkx7ls/Fm2vX
BLBJlTukPPvqkHs6L937Geasveyrc6y4b4RDyvASQCIHdW3lK4C6BEcHd34c1ccatsD2U/mEBtuI
Wj+MHrByc8xecYRif4u5rTOEJ0Q26L8IVPFLClBgzVBzUCHNZNvaF48d/zFMgIGB4Mpu3N1NSonx
0+kRC/vnTqrWrVM0yBFjVksATF+OjXIjAqxRydMd96QkE8GbG3PM0TqLOqBiwncaMrBbAcGw7tlC
aERX/8vBfMk+Nydn+eqcPW05bl8EF5TAl/EAPIKK1xV+e3ZRqlPhcA13mu/w422cGIgpSWuboK6r
frgMmEYaxn9MzAiUfb7VsUwc5NAWTv5Kt/kakeUmFqPF5X5oFDhgp9d5ZdQheE5ZvOrcFAid0a/K
Isk3E0545UHqc/wJnK0gmtxWWGtWmWu9rG3uUgt44fcTOCqIUnfOPIgFeyhxsVdbvgwL2LRBCYLd
eQuRQTiXtiXY/nHmuyscuQVntArJ8ahT/KgywhzikwwHt2pDAR3GRNYB+hsJbs8tWXYH/cHQuxMQ
XE+EgdRGrueJ/o6hkySegmoUDMRfVTTRNLPKOhjm/QDD/YVaQnOM/f/j0Osc6uSzqFTKHMjIvzgn
LT6tQpEaR2gj8o5VrIyold6qKDO0aYFI4vmmD6T+PFN99N549l704hJtHUEXeGi6XmfbzmagFOXp
eKNBTKLekaHTgbAnnXgAqNRqDnyaSdETz/1gNoHkAXMLKs+o8yqCYO7pWVgQ8svRz4N0igp1YFyV
YPYj7Jxvq8k5ZIjHEh0grVj/abBMbZvgep+r8KEbYTgDD0OjMY0sd+GXnEA7NM3M7V+xveIhhAP5
buEwUORaM1vo8ne1UThrx2EWc+6umikLF/Dm/Jt8108u6ezfF7rnLaOju5qeqNjDoIEsOE82clos
2d5HjluZ0bO136n0o6p0HM4wdXU1b2VzZlmQE5DUPU9TXhR88fYaFtDvZiryetlfVTVI1vU/QVFb
Yw9tNdZLCrW7KyfBhTlbLk5CbmX/2E7g7vq2qM9RNZKd2MCYHeSCIYSejrF9/yV/HiExqKM61ct/
27yaGgwER2xmqMTY4QWSrKvC9w2i7peK/cmyf1UMjY3gwxGkE+gFbQ03gSXTSRgGfLHfIL8f8Z16
s7NGr4HO89OZy8awQXVCmZmomjt28MbAq2GJa0N5SXJI7kH48YCF4Mdy5Tk6ImqPM6plIGGWYPbk
5wyhUUXwA2ZD7j4OicHJgH2p2DJ2aWtSoyVf1v65YJ32GR8NhAKRfrmBzeZXCTV4ffdW2SeBxnoj
ZXRGETJMZOHvPFnVv/a69YX8ae6F7H9wmUvRNX2G7cqGE/KFqj8gZwMh39We85DRkbZbutJf9YVq
HOSGYpxdl2G+lu+ynZaCoVKKgeAOS7JMFar78SHYxdnU/jrBBjoNCmCTSK2WbEH8KQhEYZVojlMh
bSO2oD8MzRJO/46rA4FMtisYoa5wk6mMD5uhHsAjPl2FMZQvofNJ/ZUQNFrfpfbrZin0AnqIx2l1
aJNGPoSGnLDJ1Oym50m6l9j4fufGoRz0Mlj57FYns4w36YOUaniVQC3tXulyeA0Vmju93BZvuyEv
9bx6nA/41x42JHOBCQLAIpGSeeH+o/RfpRe6qd4EgcKV4JmU2hvXSHtMXedqDiG931yXNUz77qqB
h9mxOxTbpLL02uGQSKfRkhdPDv6tkySVr3L1nrAnC3cRNRADttUjTNxKcpLaVbCtri5TuKhGww5a
jpqno5vPWL/b5kQRuyZ+48m+wdxU1E/SIne1Tc2JHxQECWZ3y0V413FlajvZxWRydvPDj2+OWCBk
+VNGpz5alWZ2ibizPjh5ZwrJATcI84YxbO1uM0O8r3yatil7NcINhbNAFJtHuBXH6KetTX6gxsZ2
/oqaPLjxYAh4XRxlqS3u/9u9pUjIZaCPTukN15HCzhx3Dgzy1OhBFQGi1qu+VKZf6ZPCd081CBPL
HVTbpAB/glGP0rXVxcpUf3F3Wm8sd1K/y8GCZU54+2atAWI1dO6ALfugGrNEENXoZiKfIFg5OANK
E5LMwV+05KFyuFHioovHqTOf8I4LAyEtuBBZXoIav1clSmY/dHV3FpcgH0Sda2/cMfLU+Da3PVmh
KjAjgANyDIDrQSUVjBheC3tuCSR5ED64x7VMzNepd17uXVtbUfFG1mGKWhAhO1RamJGy+5oE1Kx8
JmtKI4ASCGIWvRF/nEs4kYUblxaRWSlcnB9eTVUdMrKKqYcc9zLUFHvkZDBpxrkD5fHxsy71UFfz
UR3aUsXDEUM/N8FmElcbv74v/NNFhKE8vjAul21256TOGNSTk5SeD0OoSU7XuPjSD+p1D2dHvG96
hsJlUFjuChSn5ZD4SC8HnOoPF19E2cP8XwivpqODUbQeqNgFKi1gc2MOXqwTY1CGturXnpFcpyp2
vQwIyoErDI2x37SmjKcKxYkDRuGu73d/aBQC3PzKG+JUlczGi3L0iczQnZ19HPWG7zfiDInC4LpU
oIogjgkEevINUQL7RgNtaxjzuR8eHMEeYbU++9zKgyIGthdm3l9zY0IQvhdo59DgvEOqHlv3KT3e
A0pSbiDy0P0Zti/6dhieMr84d77CPR/iM7L/wwnwKWkdQjTpOHQsSgmAOFlRO5P9A7Gsu/4fCAdO
YuDQDFROl/Px4DUmpAKouueY/9CEHljGU8/EGz796Xm9nyJ3pw041Rhc4sxiHku+XrSCqFe7hIxS
UAGMJ+Ef3P5ULuNqrH5OSuq4NFS1oo6kYMHKVnSstI2PcybrPauR4HxgFWgqLFeTZkiQJHRkwf5F
f1E3nd5KC7G7A0JuqwGuSj32/vsphAtgwAYooR5Fcn6oMU/PjqRAVWcD0V3egIJ8HpY2OheysEA9
20lEUETBOyiR05hitSMEhzE2wvx6eFNQLKAYPs8wSUsCeX6gdG63EgobocEg7OaquwYNeIHpt6Of
qG0WW9BCB4zA8L3XL+c/zHzIxtiB0STFmLYYhtryklCW3ttMOdgY8TcZRpnOsTwHzOZh0BEQ/KGb
q7NlyI6mL98hiwtsMCoi6s71mJ5EL0ppvFT+wwFgj9cqREQE5mMYE2KDo9tOi4Y1zopeIJz31UJ2
tKRACQZGN8otpVi8SCnkLlZ74Lfd0MvWbYaXyYJm4EXPXF6bNBIJF92HeMdYgDFxcwMN02x+ZyXs
X7kG5R/p5C2IFtOf3XJx1StnFchjDaTsW+j3hrdszNVkWJBPn01FONsxjPCFVHpgkIXyGaMA1ynt
jZ7T8DAzGrtBP5E9MLY3NdzmPmFqb8LX7ynyHWgpt2uJ1pxhvPqN4SUf03ysCo394qbUaFGNKoy5
PsHBUQBlaEI3lVq8ikuOYFL/bLfaHAf+9+JCL2Qoe/94jIDYFyGD8PSfIILfy+3KjGcaJh9Y6rV9
5FWXpjuSS9bDEpwoBfdTXSDHn77ggNEhMS/Ob0i/qPZ+CfiI2VVHpmIVi108WVRgadS3ZhAw193j
RAYlYlz1J9gzE0mQniJjLiQlI4sLHBkk5HdXw9e70vnqG06JqvQgjGfxp9o0OKPghbJnLDKH6uNh
welrv+Lx5wohw5/HunqOklDyp5C0lo/NJHFt49v56wARBxEUs8XaaMWNHsy7xzUOivJyaBpuH+13
Nz1Qhx0vmQgfDE/Mh8jfYmZnMsb0I86dWEZkQcNKPhAsiKtmQSwAFedMz150RNdXbiT0OiEhz7tl
FYGjoUg2sVbG217ob7cTOfhT4Zv+kqkfTCnpQePgcTHaSIGPknixqTpLvW4ikGW7uKK1N7wjGeWB
uu28f3oXtzHtitxmlLL3xmly/FwGGFrRUMeiOV8uZAK6wPv+UInVTt1Fe13foesvvh5zLBELKNa9
Q1AS9CEc2NrnRe9gOvTvbfgRtTtpZbx1ZmAhaBXrSyfXrcf4l7P7LbCuYcqdMgJF2EIAE8w6U2PF
zJYl51lF1iUEjj5OXLWSE8QAMmMLOoW/yKoABnMOAmY2IpU18FxAzpCGXUkcxkHioqf2N5lMqWmf
PvnCzrcldSv2fmawSGHkrShbLo1Av1paKmcpH/3DCbN70iwsPp06qu+Y0IjbWgJi0qt9M2pMhTx1
B5rQG79Umb71zsKOezv61OSa/ZoV4hYFVhJ4nrk3clRHFFXcjphgZKfe2mIIgcP2RwC3iX6yr6hX
DZIFxxEYZIameiikPgnKGmen9R35wPZ+vu6loz3OtKGyADEzMLONwXExIzJ9y1KYBemYR3aaRiEd
uaTIQNDthEfp/7WyJayOOmpRjKVV7DsjBEqPoxN/UWY7CFwJYl5J/u5HRsNSY2R+nPxhBo+tXpDV
N24UTsJT/plCEaFPuuWkVhbj9PfVm0G5hAE62Qb2Kwbx8JN6nMSEwBKhl7kikHDyRDlOhSrf4T6Z
Up9RJ9iItBd9qLduQoLEEq3AnYbeYOW5qfzma2TchjqsLQP1cLy5oAU6jt6pDdIBM78It1kUOZyY
t9HNLQvnMqJK79F9RTTZqD7sp87d6reBhXB0tl0kHwJs/F9Snic8/3YIhpai/hQr5k7JaRzCSgDt
XpZNGuLMTVq+w3GGPcnsxjYnsJet6Qdkj061qCV0C51yTL9d67hwqy6c3RYRiYf8/5RNAQ4Kslcw
AvQx56DfmN7WbZk0uo4OV+TrZIaeEf/xZHGZbS4I3+p7HW07f3HRzVXvJscwJUgTyX3earhJ5o80
WMmIucISwgdHvbWEtdsUI6tE+/YRz7FkS3rtx2HSxAyhxwTa/b1GOLSotMOmHN7uRlBTNEi4CYEz
pp6vFxhp3SDrGTDevOUMqETnYNohWWSuwM8GuKvCcJihS0IHvzVlcybLCfh5WaeBnzkquHoDOzPi
QzJJYPGLEOJ47jnLojt/zTcspiIgYrg32xrPnWSebCPZrODgLunfynCWtbtJuX+efqUVVVVUhCvU
jtoeEr0VM2FwNm0TYYaU+CK4MoaPAUknJ5JdF1gysaErBxmQ7ktemoZp64KPNW+B6clDB5yKSDp3
XO71N/mKmh5s3l3sGVSgKpDN3/0DBGN8V5R/qBFf2Ss4fjT5ZNTpftdXT/WQyd+xOBYtJQY7nT2U
zRPRUDYS+o8Cxo142uqz/UaLXmOdHCG07YpnmiCdSecX1OHdn/ak0HuxAK8EvkH7U2T3AXvdrwMT
r2yqxdUPC0i/BQDhmWt+SF+4zWB0gmdh258/0S463rwxepYFAbrVyZ9Uv0mwXyIya7MqxaWoaF18
nXSVjWgXudTaAq442VAC/1ArGVKJLlJILAOdrSdO0YwSXME6j+loO79kN+5zfcCQQkIpXiOlJzES
l6KMbM/aUHtmhc4P4apWyAIyK0vSrtDOe6zBv5XVPZCQAZfr347c7mUjnzWIXhOmidPLZ8vq1Jno
/13cp+NuYbAy65rT/KeVw8vHuS8AINJ9eBCYxXSHKrEvtfRcLsWCW21SuteY4xVhtsBRR5NrjfCT
YZpIqStVPXnJlkpRVpvnIHrBNLOOlg9gsfymQTNTbvNdyiHjl+ULDCzf9oy54nn6aP/tKREdB27N
0vauEVtJ/+Hps7ow3l/DSa8Vo7v0ulCZIMwwas1a9KVJWl9U1nyWAvk2sroSgVQm6ZxwEoRE6RGm
nrPKy/STuGm3cTQtYe4aABwbylzQdYvaxTPy6ZN0zRIn9NNJtn4M7Q1V1bVcJ7nZjs9r8pg8aCI5
pk2fRJ8JYYZpzSjF0Je1JPtE2NTwm9kaOIGkwaGthDgXP8JGAWNMG6H/pmxUt7pbnykkmBLB9Jc3
sOh0Lo6IlFs4r3O8VhZPMuewLb45OPjOtXRi6697Ak/OQgeThFnNIWGsYUdoPUUTcF2y0oM6X1Bl
JNeZfY7rHHha+hJGvaSrNo4c/IsT1zHomNST5cSeON37f4WIHvW6vUdFioOwjSJMWXJMIy0Gq9XW
6OsjDMh0L3gIynftUMzfm5Q9yhP+m7KatdHMvt2o+bbkQKCBbLJGUg/2KB9qOxeub01EvXCRnkmu
jpuDjNFvg7FnELih/EU/wWd0HqZK26d9W7jiSeqXwrtvhAaieO45RXSjCFE/CJ2XFh2ysRyPj5XV
MmroKrsub8aiXqyb1Ezz/V+w2Kn3a7zdc9s5OYSFAQkojmXlU2qbt4+rwcCRaQuNelh7/AgRAZAL
twE/VF0PmAgQn7Webgc2ZzbkcO/xMjIHUtqcmsAf4kc7n7MrWDEGCeeGNr1O8qm3CC5zqSyfNc9p
3HYxOKmdgoMTaaE9CPoHtG7bTRzxW42n6h2hZ1MO58zsoltAeFNHLHERtOZlTHiuFrr7a1FPX6p8
WGjErD364ZC3JGedxVTcYLefXhVlo5zsIrT5hLAb9KHkjmnxsTrgd3EvwPBq9/ypZ1L1JPgZnZH3
H78Zpdsug851GPFEKiNkohyb3V3ZNlyyEqbvkKSCag1eZXiM4Ki+3W3CX5rbh9iOfph5vydEN39C
zLwliBcThqeK5HJ/IL/liQMf+5BAIHsRHAIetx9ogm8HPhF/g35H9+hDrGdifviCTn1BQNwl3jnX
AlA30lnMsyLE8VZE41iUJHUvkbIgz/wUJHNNii9zbqEZvF2zKDXchEMvhzUsTafAgp1zPX8FTwvt
sKIqmMAtTI/0Om95Eeas3wNle5TIQ2h1QlMUbCZnKfwHbwUKN5GNbLZcqnTti+5nXTS8yyKoYfKA
MQVvARSGMLE3DHxZOAPY8shFxbuBw1kbmoCOJTaOMslq3vLVq0VANICxPiZYT0/eFnJPKAv8SVuD
BH9GZ0AGgzUishZ2Mt4C4AKuOaJ37foCvyC7Oh/jyCGhIgeMzZCWNB4qN7oaT3cvUst2WED6UYWH
d8Z7zUdUKH58dF2IQ4NfRPyZthxtx/E97kdnnS4YyONuAbIJ0JwiMLMSV3MIFzxISXgl1gerEiEY
IcHyIiXGVqhDZbUSMoWu4218ZZ0SAKVhyQmupIuY8HEnb8BPJSsn/d49/KaYQ3DuqKa5rBfKC86C
wBMxSNcRKwqKK6Y1m/OlP4PIlHH047YkI0Ol3pDjNLM59nonm6r0zO4BsEckKMiJ+xSrbKMT6b+v
wSmZycqIZV0hKUTlKOAA68bdTLYOan1AgXwIlVuuSEOdxyk5A4zHtB3MYAZSzyd7C4dNw92mBUYb
9MBGCYW7eUOs0qWeU2eL24T2Y8D+mWRMrHazlrGX7wsJA8W8hNCJ3QtQEtQyqPnFF0M/RES3YiBK
7BZYLakHhRtfvrhncIijIngH/M2hwF8cISO70InidJOP1WXQNvqNkOf0UIv3g8G9B4yTPttaECf/
jRcfAywlfMSMJ3venL7eJUlCy80No1H9nrWA6+bw6hc3/LLoh7TOG3Wc33EcChkLa3VMgpjrzojw
GSB3j2MaEgUQI2brOHpwJ5meVXro0fK5dNcE4pHq06ALozv4M5w3JLCn7wiBoLNdt5MI+BrA3pTH
dsxHdm4gPa+cCwDxhg53Sb4BfKgeHWzGd6S1B7ui8vu26DaBm5utOoY0pgpufHgPeTCdpNPLb3ur
fOU5i1/X4CZfGZt9YAXc9cd4Q0yp7ajDQ0hk8g9rVum4To6b/aBmAWSqA3Np7EUWEDyStO334aFY
FCjEDfbT1kosuDjArAL0lCwgvLIiSbcPh0+hW6u15+kdsJ0qhGbAsnb9LhJJ6Ha2/Am93tJOEyPR
TcAG5eGHBkFYGl7EzSNNDExfbOmaxqtOx6u6ZCEqtSJWJUV4MRCdJRIVYHZaiEeKAjahBTBPl4sY
3a6vPedrwMRtxq+ifY1ulcuHnZTB4idxHN0DGxs5I/fT/QiTvHKrQIC+mNnhNihKpEUHMJt3422R
qsvpJk4aWSn6mZtiOXsi2NmHj9zsOQ5J6P7OidVZ07tEt7ITtQCsAAf4SmLRkOUKZNMfHRTgg8Gr
pqWBioxKFOEI0WMbowdtgesYg8g3kNXsA7Zw0HBGmhLUDZzlBqHF0/mx6mQKvxaP1fTXgWV5JBuw
3QkUMIH4EkvfecipOW1r3iHOmJTL8zyZ2ZsSw7XBECUi+jj8xh5S67e8WUAldzPr4I8ygRuB5QIh
Ze5MvfzH8bfWXhQVhc7ua6/79dJ43xfED2yzpn9egSwxGE4ugchidtedNQ5X7B9zV35W9MRAEgcw
tZ15esthzDzSnCq2W3d4oZgBdAwc92tx+duglB+4TaNORdHILkkSzGOyJWFd7Bt20Ga2utWn2xIC
ihTvgQyI5zjghc2hmQRaMpvEmWdjzmM8FtOBIEPBnPCWkYjijYcP0IQhEicKjk8jZIPOzy/Iowr1
U94UPzW2N//m1pA+1Ux8aaB/R8njLbCuKGS3D2TM9Q3DN9hPmTSQYosHu4ySdns73zGnDZuEBG1s
Ibqk1Qt86qAS/YyI5adG/WkV8oytE1vRVpbRexQVZOSjIb/WKa8teom2s+hSBXjdq9OyeJqO4f4Z
UZBiZNaLoLd4DKU16fYFzxgGmJFcvsLOkOj7XG0kz6SnXnlkEWZ9Ig+bIZHYZS8f9TsEVVUioVEx
Dtp6Sx0pr6hz5MYFRkAOgeAFNwf9//BD6jY8Um4j3MvJVIL2nYWzb8Hlra6NY9W5u7qO63DbQ0ZF
46ODMimRDzoP4H/W3oLvqS1uJBa6bVA0Sg5oZIiYUpXtWBBmo1mmpJVZaSnlAJkCVczGm9s8IPdp
jJrY3DEvd0wVcxFyvt6z5LlJvNxNit2yCTpy2Jfq9M/pDyGdsyQt3iBa3sSTh6+twqpyjyuR4Wq2
vE/E2JQLmIVV2pT97Lq5/7M2vm7rY9MzB/UiRaVRIRtAWOpnUdqPvAGqBja4XhbE55avi88h4QDQ
tk6TCb6n37xytUYERXm5HUf2DTJYRqZI6Z2YHXjes0G7KOx6xA+se9ZNQrh+1R75EOexemxa8U1d
/opCLCcfL5hYMgU6UQ3B09K3dMeklL+N34GFJ4klhDNhAI9eh0+Zn/k8xQReAShAhSA2ba5y9moh
+yPY2dp1UwmjNcOyIWeuG+MjdwEMqbPmLragnQuBPIpNKKPXXbWYVO2phBd0+rQ9hdQNgjkyKozy
b9nFg8Lcg2HEsYEEvo9OeNCV8GcXcNQox3PkHBnhsz/cy8e9Easqo80xq8CZLzHI6VD5ZvsizESU
gg4hz08iJF+QxOmZBjAhYDBnd4QN9qXLYNfL3I71dFP+ezw5ocsqFMo2vmr7uuI7+1XeovOlQCM/
m45QIxdA0QEC/YeLLJccPsRH0pckcn8pw69zOJRPbSdLY1t90gWeOTZRtuIDmuvcY9cluAITmX74
QvBlQ7pYBRwf52ps4wgpsQlfJOr7iauxMRwAVfmXCpBXJ8hkZ9nu4olLx2FPHJBMASPKN0zIk2BQ
KCjgfQ2fXMlv0YvzLjo82nz3hQcr1nLW8AMY4/uVOug27U6Uz9YZFyw17z2xU3OmhwZ3dQglOEBt
1oaxDSm9CjzGE6IWgzeGtgaFgePzNy7izrOfC1dYivjKEESUlw8x2Tb98WusnK1u4V6m7hTUa4ux
py0LtepYMgKs1ss9kQ9TXdFPXXRxm31cwU3/j0oQfCeMSJoFNoJMSRLnFYGlMo0ldxZAz7qYxzLw
baRiN6qszKbJmTYrFRCORWrxnNseiZ4jynKEjJj3SoLwIadC+R9uyCAuI+LzksUAQWApB5QraCVJ
QyIxifvST4WxxVwUc+Uyt8cepa1O2C17mg9Pddz5QHFd+uZ2GwaiwfbqkgT5P3AZ1q9SREaz0QN9
vgjEbh86lbfI7Dt9JO7wCSF3CjbsqO/7o1XgQL/MVzOp6UwbmKD3kzDPSuqrFGiy1Od8E4AZ68hF
Xg+Oy9R6MTrH8G83DiBs5yLqLbTyolMWUzmVsz75dSMtwvT6DiGCDLtszNmzKjYGT+UdUl71Rjyu
7tWQcHQ6d5qa0g0j1VJYiP9EnbItV2C+q6ZZndZDTIn4KHttuKCP6kRb70nQaipb59nYjZTiIcPo
vX+Dnq7WMp9L5Vjq9BiSX/A/TYl8eCvkWP0uGeGe1g05taCaWuyafaVQA3P6Y0ESdGzkW3rudOjW
K0NAOD46Qcjm+ntUusXjB+LtWta9YzJJ6friThgbEzCd9VI/EQxT9qAnU9RuQhYjXObuLVGviDbZ
pHfcbC84iouCOIjmap6x7RI70y23W9K+iTWxvhPSh7WP2mk3VngtFUUT1w+NhsaEnY2Efe8Pz8l2
DuVj2MenHcb4Uq+IYwnBhJYCx8Psv1XhECVEQW4nIKVigTpWX8+eVEiaLD0ZvhDW0nCeKb6xXVvq
I8PC8Mo9f8SkjJn/LgzdVLKEYvUrgdsa9tn/ZiBm4/PXXqubFtnvHgDWBz+LAQrz303okNYXVVIV
hrM9veT8i9dDitRMezJwKI+ZNFS2H8oqiqF507Ln9lKVzdam940REFOYtjoyiFX4d7ai9PL/fkrA
r/qwFIAP78e5DMkEaXAxwOSVha+oePJGquIHizVBC5gz7LDeUrzgOyWKHlGgcdhkDAPetXozvVEP
OdmOI0QmEW8DE4T0l5cF01gIQiKnc7dBsim7b26tWvuaN5oHH8F1KTFTvqafQQYZYmdLtb74N34E
uH6YIHgtrbarIGQ9WdfTZ6LWly7eFDua/YIuxhI0Yk3a3qq/IhtghTfnc4OdWqTUaF46zNB7tVSV
q4U5JDTw0TUZWfvRYkAGayv3r7s5WxP4lCljIXmXsPykDHJ4EZM0qqWdX+6dIL2rIiyy6WiqGJtD
YpylS+wXfvv3/+LyVrxtNb08+/GijKekl7BjP/IyAmIVBA9VEo+ZKdAIH9JEJj+Yn0imZ4P8luWj
6x9ePHxNu/KEEegJZn6D1odq9q+fpSYkbDIwJrXg6fHpQQ3okz4rSm/irArk4f1E9txaYYd9tvrh
Aqt+S3BlqB1mvKpzqk9y5ghCHpAFmypsJXYnNgqia/5Gfdf970J3fcT+r2GKnyg/1sbUF9zM/QS3
VIJGjHEbd2YYvq7WUDRxi8K1o4fW0c3Q5LuyaMq+Vf364KXJjMRj7ba8IiU6LPF8JZaWdzLgQzs4
ygvsQo2n83fZjSjwurVpyMj5yqtn55jjC6C6TGL9aQNE543CRwnIWBYIWC3YyPTxHGAsWK/FQdd+
6FJ0W0wK/UINjFIU+Bn+JSKFYZQkVX7nuobByqumtZC07jPXvTAUJZtImazf1h3EuXncbcBD+PuH
/V9oh8OcdMzG5Jv9TmelaGSIEpK8EraDb3rNQ4Ev/h6PFh/dV7WLw8PxnpORmmAoEBK/rT//6ltf
oY2pjlnpSqcu60F+qjoDJLjurH47s2ZWGdOG+udoQcE3eknRO4BjgyyvK2bdxB5xrxpnOnzsA6+y
akM/ruQtp/CVjrAjFtoo6P5rrFFcgmqU+4bscwbNWt1E0raK3wnjloxlpJ+ELWj/8eBUeSMIIe4G
Xq6BOA8DlnK2GBpHYOGLX0z8uN1rWOYOTYmNv9uyCkLOf6fC3HLvwcZYi1Vzn0osZGih/v8Yaf9k
d2S3wvkPExxwxZqHjZWfcvlM1U4dMv9IBEPVnJ/90TdQFndBGocmhZT7Da2jmty3cN10IHSPiKHM
GJVjAArW8Qy2GSLsNxzOdQ8Qvo30K/Ef0+Ld3tb0MTHt5HTVT+55eJtdvP4DTlA1Zo/i2GK8elaK
ZWcVxqZ+hccFOvHvDxJL/5ZGBXDiq6VH7txIUss9MjiKLCRQAubovHPoPlL50wfQA23iE9RYJMDe
D8pLEaVFYBqF0xRa5W2GvnD0mi2/b27f2JdTWePgzhcBsZdL1kNz04ECjF+zE9AYUxudHY9/QI5L
gl1rB6AJCq8gwVzsd7ohCCGXoWE/dsxRjcgFL3+oJgM26F5jBZSuLXgd3Zxx7yoVe1cRhmBh5pC5
ZgaHPGOvrpTtUCXH5rXlfTERwn2XBlsQYLdU+U8fmGHMDFYYGL+zRwIYEZ8CTdgHxC8pbTqnOup2
Ehw5YBK5Im3od6HjDB+kcoLq0mJPGBhRv4DtXLYRYJkGa5s/9n6itUU1H9f77+DqDSDFosHh7P+A
jUa2k77F3XLBH8eQF2j9PPKu3tSz965r2z4v64tZq2mukynP8wdUHOI42AHgqp9HngRov/OyK8Z/
fRsyDxUYibMNbvINjqEhkeOdMK2eZwjW3xNIUf0WPMHRn9DazQkpw7LNIsEtITIO6SKXRSZtS4Dy
/0q/DP7Ow/tW9mOf3+NqBmX/S5qzWMY2JQr9d+qjjhbnhsvBm/Q0YNN0foEHNWJZw5Rg6t78cq6R
eu7QPR0rM6vh8U7wj1uBxH3leeost+W6BF+aciziKMSTHxg8YiYqIgexGwhYthoSzTZnsm3qn/8W
7PPnKEhugTXV1CDrE9Oqa7AgUV/UphHbdD6VOabRp/uJ8/U+VZxHGeopBn45Bpcun0+IgQLQ8lYC
zBIb+mrQkS0lnZgKTzmRA8V2JthX/82Uq+t+FIw3f15qeM2im30OW4HBFFDK5qZxThZ6HBcEo0ki
p9qULLW+RYvlsfbueAJC572snsfwv8EDbWIPuMs1mtlVRdlJ330XQscy4Tp7TP7yTFW6iQJl/81b
wHyowAxxVTQ8aJ4KxKbMwCBEISoCrZUWT/3k8tNDqb+0g3V+ifBqTF2bHACrrPOi8s2CT7gidOOs
VuMryLWGizm1Ljxu/TfU+MB8dQ7zceSqO/yf5b1HOFJ5lN+ewW8Jfq3OwyKyobfiV9iPlC5wFMpm
YqlWnY40s+buDeNxeUfIgjeZM8WD6pP6Owfc4PbNJicIRfdrngvF8djO4ubYEsbL00etMnA8vkcC
w4A2l/wnaSrU53ALqKgKjqU4TICjv6z2PtOpTk8n8cZeQ2LjAewAj8EOF1Zf7CueqzJs8JTDgVw2
ZeMPHCDk3ypMnRRC2YmNB+iPkvXnNTBz8c5DTPedBlQPda/QAQPFQfquYde4XcAJAgSFWbnnuxYd
QTN76adkk2fjbFBmS6OhEl2hnoYYW/e2tD6m7WI4evHuVWHcjET7nyqsuP6g9+ICqoLkgtf4o2kx
C14ZjoV6RCPz85Ql5w+rxGdaMSPTOEvmCvQAQUfnubWTr9NDOBu5nT8rjtmAb+zeonmv/TvrP8nH
i9Y6NHymABTfvk3mPVXFJskQBzqHD08B0qRgEcozle13XGf0zqLoltgaDq8sO1igZgU3L3WZlLXq
GAUXXyWB4ga9IYyzShW138URjqoLdHBcQTon1OobvInVlPW2+5Fo3VCjwA4g9K6ESPwsbCzkmvEq
rhN1jBahVuB8EgIjfGhqJ8TY+r1AHT68u93m9tiHctGqQRp1MoirzMjj10Rou3qrQP1wCCchF/mm
yciDE67wTlN1VtZyElfXcQJaCW6F5FNyHx53smKBS6iUWCKBRbQxCfbY1zFruQSZkx3qhIkwO4k5
/ybNKZ/HtDimN1FEIvyVx/VHQ5fM7zSo+MlV2A5ID/CriZipZkGAz4xJDnTTSMNIyVp39DvhAb+n
h50npRs4AxinE3QzaFW0ETUz3cIXQsV7kL6S66JR3lvHxzYWkWmouTWwRPImt2O+5RSEuniW8XSN
+3J5b88N/fotxy4WeFgr/sJ93g85j1vQ9I6taOwjiHlbJ1YRvXtdIMAXxeN31jlRSE4PhW2PuQO0
TrjR1L6u+UG739Xhwrh1oOlbZnGPOOIR1Auj9AYwFVq48tODliQtNuOxhBvLtgGWy/TKyAg9gdab
1fGhKVfaUkLf+T00NSqnu/x0WcEVu4Eua/AISa6CioXpUBzThoX6szHfL83FtdKqS3o00+PDU+jk
ni1tHbQc6S/aai9xdgtZ9eAsJsSE1Ov/8eRMgYdE4NcVB9m04Rf5uf0D+65/BmLu+vH90hfv7KN3
+d7NXL9wpbMHUS1gsaB9vESVLPPYNFrwxZ5xOz6ajhk1Y24M0GwS8qwbE0LCastX4tVWafZs9hd+
8DIy2y+l7spI4eKSwwvGFmbvq2geH7l0q0RZrWJgk85ha9xZDt80aiOD+G8rYsRy0Y+zOEmhayJA
3OvgGJkQd8uZUw/zXo08s+wJeQZFWoXII2Y6e8np+dZBpPChNVR0H4zq7l8DXO2BiqjD502Q3Tan
PNTxaQdg4EItZnSMh4LBnKEAJg8Dzlr35o97BqJu45pnNnPPWEStTC1hvX+UZnV8bkaEP11JxtpU
3nwsf915ZxUARB8BiOOw8xIvGInb2HcB/uhrN8ppmlD+v3h+LnTjvEPXdXlIxQAxwn5tG2GI44a6
NClV/+bfNYBgafFgcRige/TSQdzVMEiaML464PDEL1I6aQdM5NbSp1O2BjVqdUC5x3wEThlOdpCA
4Uc3XY0T+Xa1VMhX+r5JIFEfHSGYXRiQb4kd7R2J5nM3KtEWqGb2hbNeptNxD7vA6M9vndn4Quup
Rv3hjmDa9FDKCry6AG/NW841alfOF4uqfdJqTg0TMTAHFrkOjV/HAeiOz38b08PPRfmwMtOVEnXs
P4RDxCNE3V/Suv7hAi9ufxOhdoG4sDWWqL3/8KP6ZKUdc+0AWtCX4AwEAyEn1CCh8lg1FLLDTaeL
W8RjkM9KXweQyS6H9WwnkzB+QBeinZrX1t9D8mHPlxYWZT30U1Q+UIng9hodRNcr1XwM+b3dLX3A
UgET9JL6nVZLFpRKzhl1/dNJPUu1fkSOe/GEo6Gm7Woi2kjUi32Ybvhr7fYNh5X+BvtRXfaxiMLi
Qx0n90mZg+wc6fY5NNthCeUaEryWw5f5IC/7NUBEZE05Zfu2hpeMqXEYW7pEDcvOcs9wlFdqoDGM
CRa7dIvWPZrntMqkaPZ6tM7PD0LHd5N5BKlsg+dVtZ8QSApmBfHAAfyzaJsRgRFISep7q11cWMX4
2DiTdaIYRELVcvPMCg2oVMlUZalK0cfDqal77uYBBfR5e9MvnLKaVW99dEdRy7/FU6F+QUNA0uWr
d1MPOB55UVXb8Z4LTF7RTFGaTzuQPfyHB2TCrdXcSlWFG4WJEbU+BxYJi4wmttJbUFWv6OrEMl/X
eQTUJXoe9c4Vqpj50uDv1EuVfXEZN+BeMus9OfE3O2F/uIXu1we59H6ZIAlY2Z5d9qDRZszfu9Vg
ERAHqjFskglQtcRdtihzM1zPtjzSTstsC/C9YfkGGabd6HequZzbe3+fBeDE/E8+P1v0Xe1aM6T3
3PIYT3mnOgnq+v5AdK5mXzRoTMB4y1mI5kmWyX8ZwHWmtpL8PLSdKjKIYmOBTJ6Bu9HCPEMlHRgg
IYzg5/o/gz1Zl4pEWpYVxmtcjh7GHHZT1MrqS0Ekssk7Qn5TIADvOfBqzMuAKbcCmISrkSwaCcLb
iltVqw7kfZTrjNKpCYniDCldoiVbvG9dZ9rDN7fVvSTJFY0WXLQnQnjYvf2IBgb/gBkT8F5YKL29
0UPJUFfWG8C/NKcn/iHF8RmEWbUC6OCHsUEcVXiLf87koxaXRQWUILFI5ghcY2yzh0L4gvtMal5r
QV34VAf4x+N7Env/kv125hJAbdNDLPGQ19iT4jbHlCm8G6IiOiIJt3F+W0T+ypNmhdyrYSHu9P2y
RrvzRivnzVE+4W3KUci43wG86JK0GzBAuUif4D6pBoxHoTcJf4XkFWsSJKwdTIlzwUv0s9N/HdEd
RAH+7qBP4UyLqFC1AxMzZg8BYGtFWExORTISuWccSZyiMg0qpWN6fVad/Cc8FvEKnsfDFI7PWdNq
JGWrF+c/fU/S5+UIbXwsQXIEiz7w2fOvM/xGUlhBRsRmPhrzlzJFDAfgKLgLKOJetn0wDr/KWaDz
JgZmQCddcmy5PtxBDwE5LEa0caG9w35b4dKTpRXl6i3xIawHt4DCEQyXTFFgJER4/+Vm7gLhvzv3
8TiQCjtJEajgLfAHrcni6j7EiZvKW0h/OL2K90vNTSRL3qKr7vw53d+624w6QOIRNW7NlAFPSbXl
VhlSpsLBoCIomwUhbJnPw7c5kQKdPKX+uP/fjjh1m/f8tICfOv62JHPKB02vNtt49hLo4bTHd8Nl
RYrQBKLZapbsblszCfBxPhIwD6LX1xzqSn2NkY7wtw7VOtgokWBkVUNQG979eEfYtalX5vYweuwc
9/vJavmNb4l+VaSe/rfh4lH1p296h23JIl/nvRoABcVtzV4F93ZHj2YbAAfhx1M10AIqe8fWtTUK
9m/vQLHT9QNB+KVCy87nJO1Z4Vgtb6O4pn2XSu3mcmWBVkE7+R29KhKrEApujiLDQl/oAc+j5qT2
n6C+q08zbzix/ZWzwYvHqMZ5bIDdG+RGHPrNFJjuGxOtK3sFmjtqcNV/vk+hCA42KZhsXvbANETL
uBWHBK8TLtDypIS5nvQP/gbs/j+gBO72/tRiQnAH8CM+Ba0vgX0JdfJdXXp56PJKPDCY5R3nmbsu
8WdOCkNVoPr2MT8VPVAMqLQ+y4rc7bEAaLg/vJc9fgfNF2GF40Bg3UyPu7jpXQIqYG1u9Lqnyav5
XtUkkuKrw036mlZSM7C3JBo0BiIVpTwWzCk0oUlib/izrY6Eq9Ve3GZPA3GxxcnPSG0MrJaRYcjE
X9ecqyfhre97AK6jwNSU8dA/eMMp0oEtaKL8O/HNm+WbA6EfTOOZnYaRdtmlbNMW1zQ1ryvv5DAI
KS6U7mCoFx9Sc4gbCV8hl/apj0lMK7jvS2NR+ujg8t26j4pFSr4029ehkhQ2VCTCOesH69CdRlBi
AQD0bwPMTIk9/STq9urQd+V3vvk6GFlVLe6T9d46vHQNt3tiADOtyQjqB3UpYkFDtpTtHlABgISx
Fay6WL18m1X6i6PiDxuq8AOzLVDCU8/EUt3sThfbccqA0fVWdKZ7gEYrXaAcOAbadQIjtuVzJGvx
+waXS0rZjhm3leQ6DrzSj/yAYnhNQCX4xVNBunBLzhrudCkytCo6EaXdRosARWgCFD3poCoTZN+P
BISkTrV4abdvkhXApWPZ4/OVZ/qMKL5RQ2LSt1n16EgKL35fOqeodZ0fl3VZ0RXuDjgPiZqMw6rS
hH/L0TqIf/+yTqVsoiwT1SipMbd3pjnO30hCW3C9csHalZLmFIvFCjLl4MzC4iMooqMkupw35npb
0SpHrE28wHUS+1Vv05s7KbbWUiy4TkgY1qqOIx/mRdtM2IwDPIbsKstpIwnuYMTyNzzNy2e89g2V
3kut9QjoMwBrcLpO7ZuWS7QWYWI5pS1/wMO+4frpH6MIWXdtn7s7t8d/bPxTpQAUw1UvaSY+T4Mn
Jm+nlLQLwatykoXKGUIxdAe7uQlzkw2Q0dCSa9iPWPh+fhq/5441uH4TwuOzbgTTdFqoicTi73RZ
nlSmZXE+yOCex9oNtHONTyr7jEuQrHr0e0kXNZ1c3FmBCnw8dS686F+IaV+F30wEK20f3c7URo3M
TohHnlUH/1sq9+MthEzxpwzm3jPTRLAr9+L5j3Fc7/sKjRc7c1f4hsJTcGV7Qpp5mZfW6ZpID+kb
XJvKeEqaTI8tJDpnmvUIl35ZR6U4uRKtxxC3wo59ZxWzeUrmnO4Hh55Kr4T5VHUXxYZNa/yUmxct
r2H1VulQbyfcTQ72cMkOiy4wkApPTxIvclbdsXit93Vi3bo1WLb8nE8zMYVe0P4WGKeO1yFGnvZu
XQ8izR3/97eLaPVq1rZUX2+f7Rmn2oEnlM1O2PnjB/8ICyQoRYqXeBj7kx5Pepfu/McpZm/q368t
ta/BbTXlejLJ8vvKGC9+M1LJwoDryrZcYJbfIRKva1KKqNr6jg5h/pwZxGLMfhhe/VT0rUJ5ZDLn
XflSA8KZ6uEXQEu9Imhif/jxSKRm+g5ip4MDcWw6QJnAQR8AVJu2lcCWR3qWFpX7pHUE8cbmf+2W
Kb5KdqU2mzUYuqZ+SdD/Y7mGT1wWpXoVnhlTcnppu2uNz7KJv7kGfqTQpX0MCIoB8p5lMgTJq2UN
bjttWG5j9XSazoKChzcoxf71U0E2vVjZ8RvZ5lc5cbvn/dHfjMkq6+S6eWYSlniZyvdhHcGKGYlh
Sem8EkFBqnXfdfa4KrzossA9W5oNaiyUQGqZGMLf9rFnaDTpgtJH/bZzDsfgOmLWu4dgt+a5XWvz
SiE3vB1SY0+F3tvuyhTq1dqhr9kSDiL8QAQX9xzgMNZ0KkAqEFgpm9y2Y//UXt1lOJROqLmBbhRE
5i4hwIPzEXEVonTrDc8ZlENHZvyGUedW7G6T6ZVoAU4jUikg1UHaCEmPsCioceX4SlfxjmDNaEYt
N/DeewfN7ZOeMFyr8BAw8mpKuHiwUKO4iF8E2d80n4hJnpbDDiHzfgjqJ0seE4/iC8p//WsVq2wn
Uu8IqxCRoQPqxrYWFlMju706v5ihdN15Mm23JlzGh4em1HR7PcSxXfb9nRNTyyH3Fo43XjVAhrcz
nfSgexzp0kCw4YMI4/MDc9oiSuORuwN2eBGuCAXMdb0lBEhCaWeLNMRK8bxDPIfKAuoUDVV6MYc2
C9Dm+8y2rjeoJHenreatEZzdXOoOZPY52m7pQDOQGQHEuuw5e/CLGCtOsutcASHd7kVoqSviEnSM
oUbg43fvN0MxeVI/U0mE0CKmc72tuuEMPSpupHtkTsGeK55ReJDBJ6ZPELJ7kf77e2+qdBvKpp8A
sjdaDnKMH352xtB4c10/5FiYc8nH7jcVR8eaFbQct3ixYthJ5WOv30yWeY05hZGz6K/mPLm0R687
JofcI+6blCpst9T2vkq3d6F8wnCewwYNGnjuzlZVMPKVZ/b/tuzCDSRVhg05OmGCUmOl5SRp0D7D
iftPQEieZzo9sSYhVM60GZ5c0nc2udSKEasWKOfENqlaSr4uYRAopeRPYwXVFe4fEnORK1QFBZRG
DGhn/UUHWH0ct6N5Glb4tl4QpNZc7LD7ZeiFzigE16L18Zq3mHzsrZo/+Tyg4DfAaAM1DcTWk/CN
PR1UvqTfuQcZGigvLekLgEEm8FzMVhIBnHavmILRRMpMQV7zdLd1/pn6hDLEVnaBekui3jo98P7i
uQqrSOi18T+Yy45cU9naWkMOxCkrzxBIZymtblyxPqQ2EAKSp4BZRyXOl2XA+IXldN2VO4+2w1Mc
HklOr9yDbUjxDQFo9CXm8Jf0qcY0y/NQQiCzMn6mVRvFT6F5xs5ijiyqcTbjyKmhTToGfk0Qcyeq
h0o85FKAd9muKtHXN0Y+k8CfC5jS1yH8+4c0OyDp0JmiMgu9Quz4qrvWJVOCuAfeYX7oW/sGHFjm
9EVI004bYzM0ZJDNBVGSwQBE2ewXzTZN3In4BcTk+KMQCqozPzdoxgpp+mhMKvxjH/mYLqACmX4/
X7i0/kDyKJHMWHWyvHwHy+TSOROVH0tONM03bb8FS2vqtATrdI0UUDJRYafRN9t1U6SxRqBMopXP
YMRX5E/N6HVrF/tSg1J3g4J376vypf6v933L2j+2BSVbr8guf5fxx0G2byigwdh6/lp0DzWyEeFB
U8P3i7wGR07ud5zpqm6MDVykH4mUiWSPqcYuQ6C61MXVbhrdIwOQ8BBz7ubjHLYnSYBkhuiFA2qe
7J19aZ7sDEYEcTYhFs09tCt71frG/eqcssJLL2Av9uC+S8K00c0Cxv7jlKRv65WjK2w7mbIx53gP
fAcQUk35PkSfXmDMBadcVONTsn8TZWRkLYLDCJczUl0MqIy2c45O5ELo2XLfsVC2pfgPEWDz2R7Y
mlRgdblDqsFSjMnN8iT7jRR1EhMTbK7rk6/9K4ukH8pMDG0XU1KetTngMqKb8gvhTODOaTf9PwpZ
yS17XouWFBoH5+PWkVzRPKHw+hzJ8fNKYtTcUDJfLNWSR/clNECnqdeOSDsMFxzjtoeTlYrsbLRS
WoGVyHOedJFw0scqr5Kc7PqvUMFBgKjNnxctzalaikpOAPTTnxbanYq8v0IXIVaLHCi/b21qpgYj
9AkmF/ZYc+Q8gQO0A4QAK7nvUiLCfE8J9jUCmbCvIPFUMKeLE9dqCy042M0DstXmuniTUHcHwrX0
iAKraJYr88j00H9YARoxV/3AxZaiV0CnM7+6QQRV1AowizVMDWHWSndRXD9Gmp2dB6UiWW/T5CV1
BrBIwC/8hkqgN6tXGdIBPOFerWhK05HuGNOlrYt2tMSiQP+Yz55aFCQ/oIB7lN2TuWe747r+lmve
/EQJIOtm8bsPBZ958uctdsISRPRirGnQC++K4TQIDSdTAbC5JTHp24l7nEpo0v4V4zvhb/lwVJ3N
48xU6rFCvEtOdhV9U4rzslcfugdbP3VPq+ViyjoMoRZlLT7rvrjoJvS5eEoiVPf9OqI2Rb4Zi6Fh
IQdF+4VRxWdBLMniGisp9/AJoCOf95eQTwwBmUTVu3gsxQ1FzCzwpFF4sN7bmQ2vOB02D0O0JqXf
HEL/XpAhWQV83JJaTg+/NFABXYO3ETfkQEn0VrELKHNq40crQlIrZ8hHg23P5LRXrPGD9fIneCPk
KkJymut5dRoTGj6Go4vgk06ZDJ9+xxR4fPuO1pHeIv3+U/bXDW3pc2DDELlQZlWoLCS7IC2UtSjl
p2STDnzHiPVT0n7OYaZL7Hql/z0CueVgFXuYMTaoYgHNEU4Cie/bkaoIEw6gFlW2noYXFhJMJarn
NiaOufrhEJCKJ94AJQlt/6UxL2ybTv27GgyQUBe231yE584y+ZTVXUqT2GcG6AK1oFz1c+J0Fwwn
zNmd5pVm2iBQ55I0Wpx1i/nd6lqxG82wzdY93VgwH6xOEfZ8KZ9jCU8t+hLQ6EX+pOkyVENLFbL1
QcU2Z1sfUdcm1B2SNjMf4GmQslujaxiWD5YBFSUvYYCNAa/XCl4e0XBTbMrOlVCfXELEznRs9Rk0
/c3+N9sODq39QyR4vJNbZT6Q3i8uF01tLXc9OT808qGWtsRvfydwsC5YFj/JnkU3mng8ISAcgHBY
Jhcm6SuRdQba3/DTkpG+xnPuZ960YUr7WdP3v4ur1SVgny2B1bbgR2mMi8c3Xw9wsimmAOef3HXY
uJbN4EAo69+bVcBlTxfE6x52iCd5nvzbj8nSHX7tcMrqlZgQX7mAlZOlKtMT+F+ZODxXTga8wgo0
5KUBscgOj690B2pdTUsfnQ5iSjzeREGX6OT5/ax3iwdpaDxAljrD5jDk+dUtN+OsX3RgCwtbMmJG
KZYTy0NK7qNWEKu4x9U8+Ynh8qP0Bt1Jtd1oUTEAhgrnSxFVhABeygZyuuW5Dg4YSUakZ3fI4FUh
5LmcZec0B+fbJ75leq5Fov6HxVXMxV1XSwCb6b5m4GaAeMiTnJNPXfqCFbWOLUi4WxiJDi7nC+Fp
3dKb8oSfqKpBMOpxfjS7BoO5EvcrIB8iuVvaSnqGQizMK67vJNymnv4UClUvSl+4V3o9kp9Oh1kE
VEZDo2dJotMNyMd5iWHdYloipljpv4BT5pJxqGDP30t3B0S5sNQyNNitjp3hITLarDoN05ToiIA4
MFHb682YuYtT+vt5M9v9M+RbxN0AEkxm4BrmYl8b785kuuGljXqbv4LUxbrnbDd1QbhFYCJsxTPV
I7y+SxpJeL00N9qr15uPN1/TOom13uovg8WROpebeXhU/U5t92537YihgM5l10gUjoPZiaJkB7/p
28jxqPYsd+G9PdyZOkJl2JV4jPi1PkvwbMma/MbFLM+6koo/FxycDPrNtc8wj/U9JI+DkYUmg19H
GpWGm7+OXMZOfVp5WlhGLcZXN0YKR5ZaMggo5ZNgYiDVJrBqZo5Nw3Yc2JWEc2ZKMxOJnGV7R4xs
0NZDn/0TILbVbyHy74U9eFEY+a6G0XkA99cLPOESvlamcp/4iVKRU+VFBovVi630qpiAJCnIhs2n
GUuxxzu40dyyn4hBYzBXJ4iUp+jI+7C7Y1KLINvDQkEQnZb39lf3VGqNuNIH5/CnKjoClIxLo1XW
xXXS17Yc4FO9g4BYSWMKWbyxXInPbG3iq08mtBL/cKqy6M7qR7g7oXRrJrpMUxe6XThf7jHHgXvV
21J1h2XA4tYtivRMtRIZaduiXGFZq+D6Lj2Frf6nnxmFTrMRZj4KSBPyrp8MiWioGPPqBRdTmHf1
kcUeIjiRNCqrsMYWkmGBfgMAk0gaSmB7ncy43jIOwrvPP/CNCxA9qnCJsevCQHID8k/LZbym+vGS
XbClUhy3wv88yh+s9hcQxB47MFVY9asO+4OQXLM0cN7v8PbSkisdSpE36oZClY/yJKSKCBme7n/4
WPQJrSqPDuA5RTc2hNSNIGHRJka4R+wGvj5BreA0dMOW1SG3D6Gnqs7VvQiEWLPxP9ZqZjsjfiqm
CF5hlc6Age5ATGBz17R4oQXRQJWJCNTINnxzX3ct9R6vb0gAHEGceMNjoNMqfc7jQcnd0cmQ0zk5
e3bPQN5U7x9H87nVl6gJSg85n0SBlu+RR8YT+3aaN4/241YXXZU0R32sQcpOKFOXLr9CnWGt7Z0f
qTzoZ5DVrxcwPfcLFbycH1nu56Ny9RptrMJ0EeH8pqTrNAPashqJdZYv82TNX11cZanlNRkSaTCi
zHhCBwTziFvcIvbLCM1CflYCV0qMalRqBM/o+uIY+miUue349mc/AHOFKc9CfVmUvCuZtKxlqJ+d
JqqUvTkcPW6vGU6Gn7ieZ+xDsHt7+AXl+9zJsDi1nEev6yzjwgy+hAtxJk3tvDItRzyQSFN+c/vB
kqHzNlZZf3w2ui9TpluvDRgRD3HIC6Wdm5z97wJbBfOs4/jf0AMukflqg1r5uzAkLH1PcmCbt4n5
M+6eCr3svPuy+LwefvHaxXdwN9v7h59cNUh94rOefeA6jjy2ltYCd5EpANrNy+OLDo+OvivuPgZ8
QTSfLeJwQVY6v5Pa1uFwI2LV6LXbHIVzjsa0ddAuR+QB4NvJeCNo3oOVeP1u0FaX6+APFF3ao9ZR
uIO9sRO1tCasD5vht/Ssm/GpzkCWwTQ42OK2YA5FABB3ALaqIgM4uhujLlAKhIaynWMY1SosbfMo
na/E9H5o+7ithUsgKxRqm+lHQFFtg2uxK5lso2k/GaqPch5h6g5tvP8mf6MDFaIFMVvonM0cizPC
X0a4jMPVjgxniMtHnfuoHmfRP7EAfHH/I9H4kuv1vOv57d9zg6qLa6V2gqdj5xQfOi8J261iV2NP
DOJo4tgJmU5EkoQs3OmkT33cl6DB74pIH4ViSP9qj1+KywP35kVUsEqfEhR2k3xykXTMyVgkMBLZ
vMwbX6b40tnTV2qhmKIwI03qca5cvimJQvQ/ak/3Fgk4yKEeargdoNUIRbhR5ViuVMRg97qxX+AY
gaSYyky4ELo+TNuoGvsxD2brOzzmtER+Qj7UbCujySfuU26krDdZ2+kMyZUUw3skVzQGuEdmXe7u
Jzu1PIo4Eh3FjY0MaifOaHWGPMQMUt9xF81fe9jUFUquPuDhNmqOW0EofFrwE1x4y1cFgALl+fOx
OrIvHWX1qs6v98FnZTXRceq6WhmSZnWSOzY2S6BJwQSDDgVhgF3f7744DSdDl7nwohiFV1rohQMc
OmbiyKJXir9vSXDTfbUzi2drRVeTwuwxKqxxPd9LMJX/z4AlpyeTti0mNFJjs0eV+taBTzY+/KqC
6zy8aFRPtoW6YYLQhDPlUIRGPCD4a8/Lm2SGfOg9Buwyuy7jftFeWidqxaCKM/ZBlXiu8hDqN+6I
RFgDSM6ledy2k67rTOIG/afAToDDP+aD2aa4ObyV7uzDeWzh0ITCHA+JPpMJTMl+jFYgvdP3v7mD
DtwYw9y45ObbBf64eOLPL8xEjSNAtRqsF1dEzVWA++AZ3/aWAHFtHnBeBH6EtbTY3BjmmRv46F7l
k8bXhWl1+bqMp/WA5Ad6iJmP+oty+L7VNYTawLRgI0pL0IMXt5Nn+T3ealCeSqTPcZy9+WWBtIi7
52UH8LAxu3UM/hAgSHsVCc9ylalk/JqT3ycwkDr+N1fKGkxqSP+Mb0WhOkBaStWI/NP4hQmnE7sI
43WCvpoCxfkfpsGhw9OdevREsU9TaY+qTVzs3Lyx7TwJWWmslN6SoXUpC7/Zf/HRcj31VkdM4/eF
dfZHV2ya9+kmJE3sPkP6Nkkaw1spSESMh1byoabkTsr6EmO4IGsjHJcepoRMqNS+2wSEDYmRm5Ly
sWbvcDN/+/OETtZ3C9h7c/FplRENy3tH2bTxn3La55iXMrwOBnKYtqdOY8tUcY213bTXOtVCJNcG
sMNGhGlbLXpkTJPx3dmcirHc+16c/zAdtZXCh4WVG5OeINpxuQz8JIPWKGN8NX14ESIsXlVPDdYn
B292AQIJ69QR6Sbzpail9KcfPhs/6Bz58CMrmgT8bKUZAJ28AnopZLWJIK/DcsHCMLjlKiLynVfe
HxUxR4EexSkLd38c59TKl/Z6ym/buDCc5eMOGpyR4PxAT2DVFh3rqXHJvb9bujcMIWcWNNY1Yuvs
l7HiMbh5Xg6plpnxEgoytUdQM10BE+KGljBue63kq6eebEocAztP+hEW3MxiwdQVwBHS+DMT6obb
lAQRzIcQ/s9m5q7iP055Pf5ZTD4S342y1FD/75Vb9bHOYtj6s4wKxd0BPCcqdxiE/ELd53c1UXGj
Yi9J9i/1j9vtM6wpITR6z4Pds1jEjJ+wZKHKr/4EjBnpBW2E3Kk/vKMBuuXloRvo54sJ0N1GlhhA
oLw0/DNZ8eVW2qZQSLq+MEt2LoVvor73Ac8WlKafkcJo9nV+NPRV/dZbKaFCv+suHCcQGMtKkb8p
vM2eZ1xzVooPBy809gH9nUW0m52G/m5L/8V7mm3szA14zxg8QqEkFgXf5s0LnECdNIp6oQLTk58W
dZrgcXS9svQVsojOWVAmWj9T8onq3wlaNIbCbv4GWk6Euf7WcggRlmnIIoZLGFoNO7mCqsSKOHSP
TTsNUN+ETaFjfjDd0dBwQj6PR8Mqnnvl6MHZxtJxq0yo9dysJi8SUZkmIJqOgv+Gj4c1ZjgNq4BM
bwsSzsM/mtctR2Zq4+A+dtQNPIbe8/JJ4OgZwjV7agrGKj8dLh85eozxahVJ5BgLEQiYElRiBVmJ
0/eXSj74TBWckAr4xFabXhgtAuPIm52oLYF73tMU7ZOqsT6VZR4jwE4mPyO6UtMEbGLMTrHFp2LO
Ki/O4OJfPFPjEN01CutET6h3fdCHtXXFL5IOc/S2b6gkIZRcaZr1Z5J52wjnaNQvgCmFaUOix9HL
LUBAk7ZYY6/6gqEF57flTx2kg7RowYD51eJmLYCDufgEweGcmOybS3OBem6IWSzxJrHhJTYh3CXz
C48yjBC+QyNXqWPwZZNHMMpY71zdjOwrf6BIv+BY/kOwa4aSOwL4v04fhmdvzk8zprNvm7/R4VNk
FxcvZE7K9hGh8QRY3GeP9q9+JnnFytfOqHiML1qK/A3/6DKO/zVolF0+zl182UklEhBH/e90+n3z
qnZKOxN3L7w17UKiy4idQzHCpsJYZ1rhUIeHB9pfBBna91qRi+TJSKxD5J11UNXiIXPo3T+p1d/M
1nh69xzbVcsdSwJhra91UimAdnYki2mb4QKH6xudbXM6rBfxB96WrL7SA1btgzl4yQB0nvJH0hNt
MDqhsHKwVpTdI0PJO0XJrmptvWfsqbqFjVXY+/TkBb0AcuZtw325qKuZfqBrzMEX/4NeU2LeylWU
7e9bj1B0hUQf01sQ7avex332yfyk/TdZJGUHgDZR5Ol05SpCqf1j4++nOQdgrNfUCtTtZsGsn6FU
8F1I4xM/cSPyVKY/N7FCwrVx0Hq0wjPusvLccytiQVv8B4mJLmUrWhigDyi3j9YOcOF2ypz452MJ
1iFcT5IAUPJATCHSF9nRspEDfERf9JS85KAJdta3+LDPu2YEo4Z4QMOKcRTQEONlf29syPqs4gTD
9YdmKCDdNykJzygjWHSKeDgjAbvxAcbnyv/A5oUZ1n4mwXInAYj95VcgKFV8AtI4H5V0XD2zc42q
u1p/t7MZoEXWqhwVJYVcx4ZtIU5+QSxE9jKPC/p2R3E7cSgkPaGiv1M9mk95MO35m+20pZUuD53l
Yf6w9wwEvicI8RLQBQp+CIFzxrcJoTq/r/bGtohRywd4CLwc3ezb+U4CMlmRk6mp0rqW4uqg/XKA
Um0vl+NhY0YbY707Us/PNLYmY9uUzFuWvmX4cfQlVTbCmup4wdAJxkeuK49wY42pgO2Spj11rD3P
Yg7DYG/ojHUklmVguzy2Bf0kMwl5/n1kEB7INwylQ5buNEImXwoUS/Xe8edsENIcgRLoFmOlgxDW
9ZfVDP+9UkUplcCg3q8UJKGJKcGx2zwJ2M4x7dm5oyM7YkK+/z5r2wLH44i6DGp5xyU6ain9z5YW
vGtdnduHC0ougul+niRgP0vQ5Z7WU+8TGy7xRKfsq3qu2cHK1ki2eJMyte6PopSAE9zhB8rOq4nC
KYp3RXa53vEjVYC357/SenOdF/aRSyxf8tSKbcEnN5sbwBFMq0Yg+7hJmP8wVgnqgGFfhX+nvzeP
yUWNgwiEsfhEZ/APNhP9Y8lRmfVkNWaOxLFmdRoizsMXMbLiKYtKulzGhxA0p7nK1d34iaZTIU1D
NBWaiG/06oXnB+I4uIOtaMFWtJHT1d1KfoxbU0/JW9Chy0W5X2gHtZ0AZBMZwhWgkeNipQ3jIWlx
XLa2GYHCCtl+bmhGLqoUsUd8RBpZNF8X6vVnsEUIU5Rn1slcm9v1HOlBWo32dCawd/48Uzj7DV0V
fo7L53glRYJ8mTAH9HO76vwLk1cfo8u2QPgxSAifkfEKxRY8hUpEwS1VXiWOQu69OeIoWMmqf8RG
M8eJEkXYlSl+VRibfZtYRMm1oVqtAd18BNcqPdMMu713GqO1I77/o+zrHei7Vt8DiVKaTtEKBzZy
o4pGyzJ7F+ncBf1QCXMgB1ft4cYzfOvpLVX8y5cEqf50UG5IHw7YFObPteyxZB4ukcyyLiwpXmdK
tVoFrkL4CaJf+/WqCd3Rlu1ViRmRLenL4fyplhf/IR9TK2qXu9XUIxLUI+O+GE7Zd3sboAz29QOX
OqN9tfwN9GEh9lSu0Kwo5r/CI3RynKaUpNRnSoa2It/f5sjBrn1/tjRkA+ZkItFhy4nezUK9OZyr
l/ZDNj5512AJo/PERzJROAr/tmBiwUU1ry38GBUlkM3mBa4N325m8P5Edoz3wp+fUHFcCXeM/P2r
muDFrTSDW4UpV/wckqSJb9t3Pspr87X4s99W+HQDUvjrGa7va8EvFyZH8PNECtBsn/danyefCgxU
BAHSsHF/KNXb8ktkrUHDmjo7ZwEfxJLO3B2FJ5QKMlqF2/Blquw6CS5JyVO+lr8u4BqowCA0+82D
7RF9a6F5mWEaOz56crjT70LkqTYG82PsrLF+wmAoD0DQdWYZx8C9N5UrrUL5wPuumecGRxzjOjze
FSXKyqzz0DDlrpSymZogwuxjEHTu07lQag5fLND9sr6no+uqrNs0/4rQxK7XqYLDSnS9AtDVvpK2
1m3zkcYeZKHCB6a/P3NXYWf4ZL0FcQ8bZp/BJL2vHf6+9XzYnlmCzneBvr8OuojdHigQMHlOVtsH
Uw6qsstGDh1atjdKC5+kjblBANFGIxDvKeuGow+ILVrNOb28zjuONftnD3hRwIDSo4M2rnfnBzV1
a5KnSciJmEjxBBfs4taKFrb3f7Y5dVBkdJFeAGBwhHPYHVZyhpgDhot70Tza9bPxtHN+2YjiCh3Q
YKYXpHAXglM66qbL7YW45CM+z9VQFwcCrcvzONMKYUKG4dPgJWSaqwQR53qqufYhfg2B2wEb91/C
g82PopgBy2TK2x9NGX0ugJYNIgHWoY9rzPf0hISTzB93ofZ1m7ONoupvRZF+0JserT5yMkVy++Vl
9vQ2F3ZKj6Aep1lKjKIc3uCt0uH9NPjqdoWgBg7uxdSyt0r6Md4SYAUEbvaxGNMLHCRs/jV6ViTB
/O6/8ULtmrNP+8Ztf6XUZnWs6ZtFQDAcnkWYy7KSWVO6EKicVciIXbS38f3Sg/5d+6d7tRUMu8Wi
t/ZfgOZG4KljjH2/7lnTYQSMTMUH4egHBV4U0cptcSRU7brJHDnKWwOjJVi9DCpIkkzmCYLYGnaX
Knm1AZDeVf1I5WqLreLVTd6+E104spLXQcFBw+pyUe11/A3zbDNBTHCGccI/McYxIrn4eK2f+SN/
tpNvNz/r1sO4lZrmmnnZV/6M5VYO5tWnXS4X1Si27Md23LBNJcN1l1BWlAM0ZxGh7syoc3X5OOUd
8/YGVBtJ8Yp73b1KH7uQMUTSLne4SGbrj1JLbrQ3iWPGz36dFeFbGfGjIb6qGyKW+T5qwenSEpBe
SxOsZPnkCwhupVYgCqUjijtgsEX1o6SRha7Il3O+Lfu0ywnedMXisjL1MG/FLdeIDAT2xCOVE6mV
1MsOjOZ53Fz/qGz4Dg7H1NsIJ3qgDQFV8EvfQwZ3kjtyPdYS3v7ezoeQ8kHr7xpS2MVBtQUQ1aA/
WiM3vVtKr1gRNgBpN+nWYn7yzOmHcfDeilTwThVnz1wB+VvJmSvq4sKMvGrk7hqOZc98v3lnQroh
kpV1/sTBM1EPz+xmtyrigFj/c4WPXSKXvVkZe6CJqFeDwIAgV6sB8pPbek6AenuZSlNRtTovtxzm
Pdw1XTexS4hgYjB1iJtPCYDsAQzikjZQw336wamI8OkCGGx7LfIXtMdxT0SVBCZPJyv9mIze1wG4
quTQOKtnxRcMtBNjkbbj5UhrOFmUhoUkXYX+ep/9nyAPo+uhZvgKGchQu5MGIE0nHRsx2oPotk+L
nVcB4IFpGhsodtLqGRKyJAIAJ8aqrxHPOyTlgkbQeRXQ8yUVerZ8Mch41lyn+KkUehLCgmjGhKA7
hsELocLJoDBoOsVOhEF4xOHPgs9q59rrAGjYXYfcTCaEwQBAJk/xPUVCT9Va+gNsmBWyJw6dC4Ug
Cj28ttEn3Hxuvr733vlMpLsAWQmuq1RYCTCfMqi5dasQYPgHpzeyR/+b3xSOWeAdBy+r4e+/Zg5M
WWC0ST8NGS4ofSKjQwrp6hUdJH1S8gxM0IbqkZ/UODmd69clPDzU7Q6s1ZPKK3cNn3tjppnkPi1U
rowbdUWbdxTIrk1lDJHCFaG8gn7dzQGUB32KpdJPDQFMp8is3mvBdbrjYJirH7vKv6PMqucMFYV9
nRalWwK7vbrNTAdfBisXNbk/Hbj9JTz3W+z/ShedL6mJmGQ0a6+0k5/WD5Ys7rzBfp7T+vUqOUzL
47Xz7tQri68qIkYhW1WPNBoFQmZJIjBY9lujOHy1mEtrZ2UUk7j3NCZIhE1wtHFKsvcWYvX4JDXe
gV+IhaEIhHOefgTbV2pOa8fX4k1udOknmsDzp8/GUjFC7MveQDdy6x/2afAqjdgFcvEezq7dCXbH
YR+wQHOVegIz7JGGivjB60JJGhnTi+HFIKq9EX0cQiyMlBEEbGzlWmDtXjvtpN5tCNVDbmANQ/HJ
p+O2z4E275x+lfRTtq9JX7Ww/JDo6S1G7tI0nCXm13yRUoLHqJF+nUgoYwvWID9+MadHzyi48GlH
7SB8TSSg73Vx2wjZutQOb3ARiZWfEUHKfNMhbA6XUQRI0tNP+ztYKFse1ioI4oXUshFY9rVKOl6r
gJW5Y1kzz5+2Hj0sXEFxKO7k2y0/MJ6TgEbWzis7cQiz94dBhuLO6U8H5udFqBzEHkolTgtXHWpV
qj1HqtXL9mHx2qT8oYjNBiNeP5k2LbLbFHPofD/eW1yjr6i9jdLn7vroLSGWSdhcaNMUjhJKUbO6
lRM0XpxrvMErPX+9nlKXBLTVMRX7VZhlDhNMXLqy48m8EtfTzRtb/XT2eWdosRe8rWWjeZY1frQk
bnW4H+HDEByWhLgq9GiCEGfUsAfvfMTBgCcdI/9LfTXuxCOt41VI4kDYDqpA1eYJ5CZWjXfKEGsF
6+MlrBSVKKxPao2YhLwiTh1/1WJ/bzUi0sdxhsTIj3iEH/VKQF3zgkzxpz36BEX2FvKQkGrsxYfU
74+aBREBPBvWRfYjuvl0Tp4UiMDeJi54Gl5IYrUsBkLpLcDZPuPR1nxCDOj5neeK40m/i/PRjFec
QAAHNckuYQPQxErqnqeojsxdzkxea/QhiqrIRvN7y3UZ1FuaHbTWgnNo+m7f6HsLZ+3CrINNusm9
GDZIauloAK2CJUbhDnUVBF7Fv7S/5hg2QyIb6sAM4UxdM3FjeXi6ugiqa4fS6C/P73Ggx6JOfsrl
qElBGeE4407nUuqnToHUiNvPpstWI24OxqQMf6oOzHjkuiyVaA1mAohI/q8/K3JfhUBD3gL8BowS
h/Hiv+Ymw4yML4AX/FSTOZAt+AYYB62laNNMTgYw9oRmdFOMWZP30GU329SISJs/k954AGcdv4mA
ulg3f/8QT/BUznQh4hllgz395pa5jNK7xxTtdz0cCBmM4zDUn+HR/y5eR+V9HI8OnxHXiVsoTR74
L+RbM/DHTR1LY6bc49cEwsub0Fr+AzpyYySbM6DBT5hxLCZ7Ool7ujqIo53fvJ3lUGQtXR9dccOE
JxOe//PrRg+pm7kwzsDdZzOAlJu08EajIv/RmrYf4eGjbtkObpRqV9u5t4ecXk9++LfBQXsvN8M5
ZM2tEWNCUuQiM72dnUOW3i0aVbv8MzavY0X8twEQYpEA2+ZwqisrfIvMNsI3oKxfAKs8QR8ibNdQ
qxMBfZjM+6lYBIHth4bOCFqKm5aTsLiW9QWg4hxwfJ+a1dZVQR9bGV4NmZHx9LbRPfRMfJnQ+7x+
bcWrsEbI+k+wNTexubHTEtAoBSUh263NjgDsVDFJXVcKz0RAKaFF7n+J5cHMw9GsR6ex1mvCxc+4
82QRoxzUoF2VMMSumZFTXdb/cTtEIRUX2oFxO+/071g5CNOBgfyw258fykiJXDRKKh27sUl3xUkX
N9kVo7G5veQmSR3YCjJ1C4eV7eNRcEUVbfrg7E/+ulaSTrAk94DBvRAC+w75F/LDZmgE5iFBXLd2
Lfs0ONU7PjKHytFfSVsVPwDyEgpSOTXXAaXKyAlVpIdGKNRVSS/2Tm6S4v4yhoqaNyv7Cw91Sflr
djBpkpCiw00oNfhHvwTBry2nY1rEgBhWLAAPeRamAM+R+Mo4/5I2qb29vY9s/iGNNJy3Gmeafqoo
/0oyW1RxMP7fIcOiZ8HZqn7RxAvhF+JU44gXi6cd2CbhdITV1vd44uGXj9GtvuduDNrWnbwMMZbQ
BKQx42OTthxrK41Rcnhz6GQTxxKYRQ85ZFgFkIDi/N+hpEQS+HTdfQV0b+mJ8FG9kwhKejlF864u
3yhGlqpCT1pdgrZf9cx1YZnSInDuW0qxlaj+EwMPkawRPwkkxS5Ox/r2QN4tXYucHVjEo6mH/Lc/
lM/Wl9KRYpyroprQ/xrR6Rv4wlW+F1SsFUOLpf46wQ2cCpdndIDM8FDVAlr2ReI8kfPawgMl0SMk
tDJeuYvHgx51eLIvUFoiStE5dMOHQeCEvIS325kVz5rt/ac8nucabk2QPLR5B1neYFER8kWMUaRp
TxLlfHj+lnGk/Lwr/c/YtvMPX7URd9kjsYXJqQhj1qPE4LSxhXfDjutpu5ujHwrv2M8X1KV90P/W
kT7V9KrCRq9gb2xnoRtjJ1J5xblPcTHeGUs6HrNHVJygOWwYaDE04zMLS2AnOpSNGuVuSRfxryY0
LyJIQepfkakW1BfmjP3gxaHnE7ANCtFENf7KNpI7UaguJS1MpGQpG+lOtrTDXiGBzC+OMgSzHN40
VVLhqG8PDv3VR6etIyCQWNpohjCj5bulyWxWKcUJVvIrV5lLuhHu91C7odFwJXDmq7JU+qG1ifoY
Q4m4R2sncAl5z0soVdcuRR/kkcwQu1CnZc8WY+x4GlPX/GwUB8UTnFABmdobYTmQqHQKXZ5YDfJm
QNab37IarS9xqSmUk2LSFf6IgT+b+ZySN8WWuI4kOSA8QijW2/a9418ZK4fG39kJsCmg5qbddKla
+cUq7WH/QAGGr5gnnrpxxFNpA5BHrxYJ4Y0n7Q3Hmll9oKoNISK/BC+7T74XS25VSpE+KtKXjGRZ
oyNKnpz6RKrwRl7SaqgCFoAqK6ViYUqgNdsAOO4Da/OB1tkUKLk64lGAnFe6YrFRBFrKgQHdp4Al
6Wnbc3J9HjNYtfy+ixrBVD9wNm3G5SedUJbGU8Y7Yvm47yRx6BhAuCOfVI+LhgsmXfbAH7HPmZue
mtmPI1KGvgOe2AN9BdMyMiZB56eXiw7okeGNg1kr+GSHu3jaxnQNPifDqZMG2twjsTtpkWSdksW6
mQfNWQPOSG31Syb4W78/50pcYRjQUYj6Oxnyl92FTRM9U1RKlpHYx67mn/XEWoTWjd54k7SeSBY0
Pm5mvTt+GYcEzsrGkmHHkqLhL0uA37usxC5TMzD34ONG78RjugpaIZk9x1Vrds6aMhuPmwe3/Xo6
nev9NDFEU55vZQEPHs3NbKPnZjQ1ximMXY0WP0WF8m7QH5tAa9qhsLFJybJx7SIhWEU+GxSiPk9r
gsNxDTmAzOBMDpYX+aTMlZR4TkHets4wqeoeJ/cRoccZVUCU9wqs5XTzbQXaiNV3rhyU7gmbQkls
4FQEx81NFUWEcwNhuVfO4MGJr68HA5Rio1cMP++pHzV2n8YJaW5L/BzhxkG9K1EkQi/DlFWzv+NE
HKDlcBd0OPsoH+bsaohwpfDl0VJdNg1RLFjDp0vDhKxQv93mpDTlaXHlONTKP30tP58cFgGP5sxA
1kvq88RXYPv1ehvnAQqUHsW60bbYulQfCypa03eEYkxBbVOoTXJvu1kwUg487AIHenjowNSJSHeE
/JvzSbRJkZpY0Cx2nEMEFYLG8iWBaZWq7wZFJ4rx4b3klkzknk79nHTjePyQ4F+c/kADGpFDFgjA
AvG+ewGA9Ixf87LA9BuaDftb7YSqIZshUM0vLIj6x+Aj0GAxrE/S2OuS3SzyQuQzHGCRjU33GiAx
VDSdOwrEwjXi9GlwC0/h0y56NtMBMWZDJ3Eim5jl9aaYtaC3GlO20cf4idpHXhjT0ePfhg6KeIKG
9aOQRd4nYsEZdiynKul84/A5UCHTq/8otCXOwlnSRu1vDHGZmwmDakKnKmnfsA5nrZXEJo4pXrlb
PVBzmQa+UhASzb+o4OOauEVxqOWY19VYMnUZ/cqPPPsT70EQsOdJHGAAsernsmFgj4y0XWxGK9vW
t234gvttr0TuFAv49lc12lXlHdQDyQzN0Wjj3aYfoHG8YfgoC6PcS5Z+RA216dUWBayIuRXt48q2
A478WY/kjCGtn2I8TUieBYJeW2c2Uq/u8ufvZ3b+gMD+lOQP3k/b5TdMPXmVr2veC2BuZNas8Xug
sSRZw6m6yO7kDbPW5b22byr/4BXAY2iBvJHofbd8HnngOsGPkdlF2HMXJK08UzIMEaYpFV9PNytv
ORjr+6+wHw9K4uefo+PE7fTkXSoy3iwLtMI7HG0UKxFYaJQudzMLNmIIn+nkimEPU3XWfsSRPh69
oSzFtHFgZPyvjQnHvJ3tkxBtpvkcmyPr3lnm5ycBp0fR5mEtrL9bSExZ3J+eVZaGnVbFBTvTZz0n
75N72dQ+moiPof148c9F95HyN9f2CysDDH0Mq9hFmygjL/8XY+YgViXu7s25ZkL+gj07lFNW3Klp
SLdTg5Yf6qOrL65K5ggd2489WWfCFo61vYnElyQTP5a9fYr4c2zRRUHxXAbw0kXyjruXPoOa0z7X
V9Bo5zGrhtFoFyLMdTglxuWGNAfmU09kPccjj3DeOqIs57hcg6gp3uPgzakjpzojsKMT/7sE6pzq
u3jG+YXtqLoGhG3dKK3m4dAkHdgjJYt1PrupaiueelnOR38k3KLvKJ95v+XP+vxYNMMn1/Ag/0qa
/g0lYmurN7d5npk2S4TgxM1Dd/fZ/D+huFyjf2+885MJNepdKQaW0jMWYxGC/2H3wLaWG+i5gRhR
ad2KioWjriy+0PPo07r6gMWJUsZCS7GaprcgEYC4jD6uyOENT+Y2iYr6Iulu8pLGzovAhWlc2tdM
E6S7N3bJp/omO/FO8p+GPIsK/hMlzahz895dSLYT/tSI6FHVEMPD4q5GbBoduu+Efgcnc5qRGGw8
/5dhhOaQEEcCDby3Iu2H9FftoFNGxjwJJZ/7JGucxEzVy2CoRAlIJj/fYag4mrhdb7pqsX1eBLCG
uo4Ro8XbCqU+xgNkHo9dBkK5vR7sH7Qf0bkO9QO19qqHdjG6Knea9I50XeMtImzmnPRrd2PyLOQ1
C4Q8DMN0UfQ+tssRahunGFAb3uRjFFa/ygEtvwRyt7O7yBI5T5X6bh0UwEReHCd30tuW1GkqiVF6
sYRqPQX498otQbljBPU1ytXajyG4w3Xu4gMOjTJekqlqIlLhn9SA3ztJ5ln405iR/J8wKmYEHvCx
kN2lSp+A7xYQS4+/Z9EFfZo5errmO45JXASx5WrgR3x5UMosAPIQ+P+8YbgpyryzBdU2q4LMtEhR
GWEYxgi1g6PFfh36QXG41kUXQqJE/jf7Ioof7JPDPaUET2McWgBfuWvgwwf3YKdwqkZMf3MGmG5u
USeJEdEsfeHrNkcEheTlzsOIgGWkLAoUMgeaZEmYgY4m/AjDdwThdsamvatQgLLmtkMrFFrRkJki
DCtKTm3N6ATdCPDVTSJrR4Bh1nc732SMNHkiB5ePCSyb93Ale6dl9daX4ZSvQrpx3kQinE95Ghuv
6qj+4JF9IbRFYJS6mZSFg0yAShUtvfqS4vwvUF7VqRUK1xAtGM6P9Bl5V24ZcvKyMyslNuXg1R3j
FXjopQrszLOE0y+8D55bdxBxkAkkXHoEENiUHBgQDJwPyVz7pEvwJP9t9AT7lXHIJGTGgJgeFGvb
1LBPv46CZGIwUC2lLQrhCxjmBKUl7cfKCpvha2pVUPjVHQXKDb8FXFcUDOdkh5LgJkuegLwYeFU5
bK3z3ErjbbevoUKy7CkJ5oU4pcEG2aUH8WlzjlH6lKTWq9aXTmfcLxcJnfnjVE9xBgSMrnlxnu+k
tvSCAQ2XvrGJHoJ6hO/HaLU6QV2bboyl8Y4MRTMP3Ss8fCNp1rKi301JPE5Pag4XxPNVxCKRsqkz
CnCRINpMwLs+SXzf07VRzDivUfTNaMOYHAwaAH0GSvHInE7gQv6rJCTPL9G5fh8hR8kbJQAwQ4+c
ZRlvlJI6Ic7scZKQXVk/Qt6xlykkwi4zyEaqFqWrOU3+BiJyFPKb83+Fo9/YOZsqzt8iJyagMsmf
SGUQRqWul47TomC01+rOdu01JINKc+MRaZpyDnQzfu2HPjnkPJQ8AG6THThT89xV+Wg7/4FqJ6ZN
UaW25pDm98k4+dqltUCz8wzFH+FAcZMxzW6k0Nziy9hYE2V39YLtDEFzRkDijy2d8uPfBGUKUQg+
C6MMCvCGQ/xvk15sF6iFUSufxgdxdweE/ixzumKS7ToUQmaHs2AEPiGxQXTEeJY1m0Z0oWpazbce
Bl0ABY6U5d7nBynHGk0pCQ09D0BQVanPUC5YKpX1dhNPBmYKXNTl8gBEYF5sUDtEvDYKFye3xfKw
/DE22wsE/8F8zOJx7HU75TfJ1UbttI6Jf931JApFX6OXfLfFsdsdAhl2Qim/XCppFiv24nPVoPfG
WysSyq14S8amVslv9aVPw0hD2JeE/9g8yOnrnnay1olGnZfZXXZUiyx4FEgZbZLkKHp4S2xcYbQz
De+5cR3czQr5DXf0WzooPtqIM8RyHge2HbPdxUkEgQ2c8Pl0q+jV79mnwuQwNBL8tF5gJKXeUrvq
UW3gIDdW2wxobwzEvdC+q3O+tuzpuTtxZgFX5abpI8E2jECmv+JVHbzLkv8NSwwF+z7P0Z+ozioN
S8oXuEH/VksTgRU0oSAYwYeCNnig/mtryujCThYjtBP2ouXTmX2Y8fbx+X7sva0tKEkuuJjQJWK+
ngqnrHszJFiOb3Y0yGtFvZmaQ6fjDj5DudUDzhrNrqYbp1l3JQYzCMIXuc7/YrTs0RNN7NCdjpp0
XldDCQX/fQOsLWntft2+RfpWwOPqFzGBYhCfK3I1NIaprkgUdHMIdCfpdH4zk9Kvm7sONb5OwIBX
uMWZDv5YELza5hT/Km80SbzbTnprlHzg3Sfu5gFAfxQlrqxHd35ALZvt8Y64nEex/J7YjtkBZMFE
X9FUmUJdxwZqz9J50eBTQjLy5s4cBCCmrt6Sdf/WAFq1aWDEaBJFR6EHStJ34o80Yqd8pa/S+qQR
Sc+4tdznFh2MixUzI4yG0kp3e8r8TYH7lrCPx7OX9lc0L0xcM0mtLMVOlhnUx0de+osvUU+cErvF
Rh4WExF35Npkt8NSDnQXDEenjSi81eq6LVh4yZKhhrFJoROUtjuxnHyzp6gj3DISDJEQ+uvnE2bf
dIHjO6vktxqXGaNpXzXv046JtcIgA9iYdPmbv6Imy6+dhWWRlkPF897Et2LbKTDXWEosPvQOwACn
VALT5x5pmPkaaMLdaKESmQsfU8781P3L6Afbbc8dONBniMzjb9YU7rYTPkBUUBY5Yis+YTm66nsm
PQLkvZUEZkyHFdxAz/Pc4KNP+Yebeorr383G6BdRk/fo4ZXoR4RF/2nR4UBhCvdKNNHACMUe14Pb
tKg/dDq9PO//41vzeakB7MLIk4sOnL8C+yicL3/aG5k5yroGvagaBP6U8/2tAKFVeQoTVTzU1o1b
MHDvIvCeDqmnP1pSJUXyNFaX+P4PYBjBtZx5kt/+LRhA9fmW7dygwnSVgJNw1OcU34dVi/VPx+3p
eB4liKJv4tv6lklWSbkg9Ls8fOYIHOxPSqmSv/9+gqS5Fwar17XzhzWAzYsLWbrONSi1TEB1+7Hk
c/1fAdHgBpV0fZ3MAe9t6QOQJNRBztiPLeDqxQlvCZkdp1b/hdubwVTnw0GbEHGyOPoEdmu62GwE
pV88ptGS+KMNnTmwB0wO7GmNh1A2ToAsv0pAZeCoLW/TinLZycCgwl7ulozbpuGxBxJWj2RaRsyY
rYvKmw8nZIn/1B4FioMujph8wOqzmZ0el6BjQCNPgCRRQOFj6rhSASm0vlHupvQWZtEyex4dm74D
4G1c13ZVnb/4deATbya+18hgexcQ+AxXFrVG48pXNdkbDwdiDI7ol48plig0hmACwMVsCBW43Q+v
afjQv5WyWRwLRuRV4EowBWAfCBAVv3jWlNI074u1AMBOgD8qyh9ogqsbm/I11kMm8l/+ScYI8NXK
/u4ncFL4O5VlAXtPihDvx21IiiPO40c+LAnD7jW+JD20XVhvibDwRHUbQUOtB6LzXodzz/EZS0Qx
0SsB6UPnTKIJDLe2bCI5h7N7z22vwVYCkBapBN3/17uhxEy7AeAfxNa9GAwIY2nVoXnOWSC8JrA7
hHsO/htBpcQtggNwAgRT8LnhBBsvvkaXy3LQ96OY4JyqjIZmNzw0GD5TtDths1i6ScFHZEsULrk6
DfEBJDbbjUB17Un28qeZKN7/nW63HYIjhXmNjoVslFRNCLYK1G5ysXsrwfUNer4jDI8eQ/KZfGNN
L9IiqtUZ65Pc7BZRRaysl30eRHU+9BaEaszCoxJUO9mLUk+j1C8pLuBO3UHWcsm2VymV7F995VOv
6kH40s377Yqy6H8Z5lPjG4cz+fgB+qU+uSRV8YZn375n/n1s80Pbk1nBQN95A43WAAHbpTLel++/
S7Key+29M04J8A9w5nfFhUHu/vj0ZFetYwUhZ0zTFvs9E1ttYWodRMt2lnEI+TsPaXW5NMHoCIjU
bxvTQWQN9X6zvWveLvrta0xpnBnfCZrGh5aJN4RKgCxOvzctljfiW4NrYpGlzgh0T705/imQsbJe
rYnZUhcsGsq2g7LFpV/NIAqJzNjdGBf8FLn1lR6ZxYS0g/C8TwLjWhMujwbi5q15WwVHwKbyBFHU
r6rKUDw+GOBBSSK9FtDLiVARqZgOc5pGn6e5fjnc1PrkK6/IUhNOq8mQdf15rDRKeSS9yzt13eKK
mRfNh7eQKWQ3QG63LoUCj4+vmlQRFWs/kxy8eOcVyHP3ZPwLIYnJWOf8aW5dY6jTbnPKWkYbmCkw
q+qUaFHrdySXyFaph+4+myR41uLjcV+p4XfHqKnJL8fHspq+n2UspLUnN3/rMaWvRWwL18ZuPScj
YKBfJyLfOiR+aK8ytljX2w+yNsZam1uhQLcWYlbut4OUL6Lfn2BMb+GoE8Sm8s3pkwDFBMXPgJuD
bqbgrPvVNdrIHgNk5ZEdMWAyAjiLEnWB4Mz/jXIsL77Fwmik/kc+qBtAmiuV2RJvxCibSN/RDqJ+
8IfW2NWC9+GKknriq/smfrJ3/OaH80yysxpxhJ3u96ZQEGwrG62cEBcuUwznZ91LxntZXoxjr0B7
y2VzuVfxNcSh0NgWPROP7thWT31e44UmrAvAuCgloHA6laIzj9BiaOj7bvzaLVKchN5WrQpWoHVw
MaatVyEpglvKmryj066cjpvl2mnif4rdDt8kb8JZkyso1+CGOJtXBrz/Zu/HvPajiSyq2R+YZmla
FjgP9VBvEN+xjDYgfqeyGveyenyp9MS2fvX7oC8HpHmtTFbvtGaoN/RFzqJZJ6y1fBXn8T4s/W0a
lGp0qOak+t/9osSG2cxq29zuZ9d1Jf6y7zu/5D4MvYi+73JRX1xn8p9ZW3ixQ71Xl/chBDGgaHle
bhA9FYFUJWtx3fYmxgDq1faU12s1+viBk2//VUdcst74tDH3n6Ko4bz4+rzpfb1XfrUa9u4hJfKy
q+ECJuL8g+f7vEBApRVtMIrjH1nN3tINLEWZFBNPkdLJRirxljCVvH50PHGe6AUkpBlsoGBUoVI2
KX5SbAL80XWDL6E/63seP/48tQDoFatal6WOThNUfvLwpKg4Rf6+19c86YOezNusi0gZIK9gGn8L
KKZ4FDYTPBURqXg+0AYRHnvGntD9SYmDo5YwkGTTknWuDhWYEOmVBKizUOcWJ1TicSBpfDpaCpdJ
73tZ9whOq4fhSyNIjrsqBxa7h0Wn9lgpw/vbu59viMHd4KsPukx5Ovh+vOA6ZeqdhvF1tPHO3GTO
L8DeJAnaoe+Lez9KWpxTQHcA0oP6oonZmc6v5NXf1HhuJ64ofjdqJx91QooByI6lslDT+mWQa+tR
GAxwuUNNIS69poFLPj2zAQ11DrMLehAhjiSeaX0Z4uoG08uCMGNG/1dxtwET8p5w4BPMijfIxrc+
qhJi6fr7ntmspjMZm4kqZRDGEBDyT4T5uZvxtmmWymGHssgud+HY/7Ci5scM/+5QsimlIJygPQ9S
pskJs5yzdQOWBeCIOrX1pTYBaJK4Jk1GsiWkUhU7FCwkQgwD8u5TbOJq9DEO5YsGuTbLNS0CMAnN
Mf1f5Y1mI0lLP6ymp/K8QVTaVssMOl/+dPFcwNv5jsF7SMtDxUifqnh5WRvxnxaqpoMgbMDjS498
Sc1fp9xHu9fBAbYWzk/3WLYJsq5DQhUURrjoOE+nxaYZJI9O76pz0MnApEMLTbLQaSJL1VSJ6ri/
GMSPqTNieEsE2xJLAyCroBNLTrDvLJDihHi9QxIKRpO3GEmBr7lJARto3Axat/rowQbWKqMhNm/U
7/BgSFPAXIf+yscf3ITi4GmsZXQCnEWICU8bYtiHjDdT5vXWMsO6qZcZcr/7RvTgiRULXD22+B3/
juMeUrQ8RUU9JwySV3lUiaekQh8PlP0G871jhgdrN+u3RLEcoTyp+mDi+g6ulDvsGo6wFS4fPBWM
1aEkDPVV17CepPqym+FVJx2TWAxbxWef4KgkJK0MbSdPtavvjX7SFvs+z0Q0E32MLmIPO4GB60jp
aqfAQpTVRpH2sbjwQO6c5A4Mkt0xyFFKx+qlGIq8gjEZGsRF6n6eLXnhpKSwgN9L+QpANq6W4PbI
llaQu9JemefxDHzBmmZvJV6KJI7EVJnr+zBkzpk53UCs3tC6jdeHcCf1zMh3BCO2RpinG+nxMXAr
2DlUJkUTglDMStMBBJ/MJMlnGn6qIDCsYe0xO2UQHCNR1KY7PQgwPhg+mr3eSjxS6XhKsHqzSuV8
va3B99kYw/sLxUpsmev3QXyoiKqPoG+QlNF5GY8U33Hrg0p3JGu7ClxsS5pUnMq0Y10sRoCZQrFY
e+Hr8Hc5i9EIlScWzJmJTR5tvpB+wj1BTvnX0og79LBsDwUurSa8xEyiIpWUslz8wjgo+7vyIUJ/
nEPEZUJYCV6W1W3nxKZ2ow5DE3FqS6GWMcTdjKfQpJj3kaaIX4y62vBQxvrHAdIxFdzlpPYjEnN8
M5rO7fzaC/Od66+kwuw87ncKlyevs48J+feQCQXc50dObePA8mCKnRIkCAyYG0Zn0HPOmjoIFMza
lbbaXSW3GD+3T/DXmapI0Rx67vcsqxUrsNWqaLujS27vAIQb8xtC0/iHvg7/z/M3bPxbEQc9f6VL
rRJrO9lJJzIByrQ723QIJmKSmapicT7a83sD8d1YFld+EPSoXdAf6pkq6Vb6tVLcVZdHsVWzeq9r
X9Fx2Nau+yKUvmRbIw9z3BatdSVER4RPxncXDat+AXxGLKFmE1RKnJ11JANAppZbc8w9yiFx8zNe
oDRV3x852YBt5RPx1AW6qhvTdH18DtGRfGqBUDDP9jzmoER1wYkqHSbX3J2XXJUegiSD3kG+nhAD
EAyNthzhAolukWx1TjVaE6P69EXkXc1d/DCqHriQwKEb7Zg+ylF5F/XTI9ip9JDCfxr56FltUcI3
t7pWdaz57TPDvU5+mD5PVamazKygQ7HURQHUhLfNtsbT82UJzQvJqWJypeLx1fpMVjTUa3fhX0u9
KKyfC2NXNVvA79mbibgXiTqxLqIpXprlkj9VCApmTHN3FHZgTgS31vQ7XosE+YS3MXsdPuW+FPhT
eM63GfajGjlZ2mtJ/dB+tAXUer7SYLpfOZuqwjPw7ms7I0OC75iU360BQsYDj+iNtlY1rUUlFi82
sUXegEmEVfSh7PD3J8Cdy07F55V0h+Bjny4DYNUb9ITbLPvdgZ+EQidHlhTtGmL3TzpJ3DPwjfqg
2NIW9kKtNnYuHWQN5BQusew3vgXLnE850P/Sz7gup3ULVXjvuHHDYHlexqIlLGpnUnqU+9QSCUUe
BOetT+uIH9im37bOkxaf4ihu0/9dj+esc1mulLKEUgESSNUPzmjdqKe5M7Rt3sHQaSYXUgTIGk99
3MIjrCvkWfxRqjCqxZ4qZNFhIKPTE5kj+JqVzeqQGJQpEPHx+AJXnNz90M19hL8FiiAQS/oD7pXK
lED5mZgfqSJvT5bT6BPV2RwJjq1BysKKY74Mbw2n5qmzBNUk2t4gxjiHEHB3Wc0gw6xsemzVgAOQ
JF2sXUTAVEBEkxBBmHw1QP7YpjEf8QU0QSqR2dK0rfjguoi5UQd1KT1GsaV5cb38TWf5p0NDJg7L
lx9m2X9m/GIbCScYQgTYU5rjqOj5iYYm/nbey6w4Uz7n+mwr/sbK36hDBZS3xCrTKqOWRbgPaEas
qpgmKHuVfFYpdeF3lzFrGn4HE/WDw69idwIzLZB7Jrm4ltawinFQjd3yhquR5GH3wD7bAgkc5Z05
2jt+r0v4v2q7Oh44M4KbsXjKgie9XL54IkOCl/EpJAbkDdaPrL9M2bSdEOJFTzwoWuHOPvssk28G
I2vwoEO2ZtcUPSK3rR3942Fg3ZgYmzsHCq+LT6sMNfANIr4Dan3clpkNVUU4Am3VIQPCfreqNV+T
mY/w3G8163cMpLu7hKooDY/bwsbiRJ7uQlv1QR0UviFM4iHByx6DWfzgkd7cFjnEGfDwV+HMVXnO
wymutr9tJYB15xemU5n31hDYeE7tdUmxK83padNRst5PJ6K/ILvISHM7GbGR8dAQsR7+jfcm+lSk
7xssbiTeQsnMccf5ZqQRKMRXtxedv4sZ6SQrTBErii6j3h53Hq0ujDkk7WmQA0a/MAHArZt28XF1
okHsGOhSiADqEx77Wc9Gj/DE1mgeZdtBThBDNOtrahFFXMFuis67jKKu6hfaVkbTVy+G7bywKk7n
9PIWZ5LeJURg4yOGz1AmbWCiVI+HCwm3myaYE5/3eKg9yMPVA7wAYS88rtCUX2bys8kOWabB10bv
DOSHHzrbncP7KXH+oKUaL+AHdpZRd11fFWb+/Fa3VZUXK/kzSkqnJVohfYX3kQ/y2NbLPKB8vuXz
rDpQW5ssxOQDUhTjEPRn5rG3XWYiVOrjSZty96In90DtNHf3nxxEGB/F5a8JSf9B3wbOSuT2BWGU
j34MOmWULJIFfLzLn9f5rIKvwYiFp44U6pfkApcdkokWLXQS+woVBWdcb6ySxa60WOyeQgp2hZuR
p3zP+1v17aEfZW3EUJWqlgV2Zw35OKWEOPYITuth5YX9emMW435z6Dx3jCwAbQ6RKjNRDWN9wJ0c
QDGP8Zb+C77vtGbOCyWKYKBCs20/vGIbOz93bMZP2MSSIJ67t62bEzINu+1uPD6AjS2/A34lsGLT
omdcAWSBenxGAd+zTeT34rV1sHni5Vb62CPHJZeRYnEAlgY6E6tlBY1TvCrVKvPBf9FSqik560Ww
ttbSxA1g2vj4sNgLtO0DFl2AIi0xmokSY8LOcrFt8cUxbB4R9JzJTh043NdGxe+CBs7n6hp9GJXd
0tMpsYmAR1AAZtkNmL17lfCrBLwNDwCuRo/3+eoZ5DoRmpVQ7uPBMjvcLGKWcL6llLN9uB87easo
BHx82LQIJj79m4I1BP6jdaVMGTBxEXcZBsCEywZCK4UFrkYIaT6uM+yrFRqhEGYGRbR0iMkWJuNV
9wKNQaBeZNMTmYUKk37CH3gNlCXDSm5rM77xIKn7+5+P7atsL6ex7h+lteXPwPS8BtnIKuIa7ab9
BfniSKn2XB3nN6L80bb4alBEJwE/6tY1TIOfbeMVU8crZtiZV5m7UTtC8XND5VrA7+kwx9V5eG8L
wcxcFa+8CsdHZYjbS5QiLVuekZ7xR1EissXT2dkxx2m1v8AWmo/gtel5CbL4trsnYc+ITpLjpnJD
sI6VzI1vp0PoWx5aZclJs1NFh7AI9M/rRFYaSxKQ7i2JvurrcqO1irBGxJI1HfQc5SgeVjJDw2PD
xHg+Swn7OenRzK2nBaGE16oNCSYnlrt/qfAAm2eE9EMkBi5BxsIjA3Umg+y25fQUvQZc+aIQaQ5n
sjZD27AvBnwlR39hihc8ObI+IaUoEnC4/MGT6/RmHWTlW4nQdTaHP5q2fapc7BR3a0AncV/yzQZr
s33hnTs9W3XXgI7nsMnJr5JsLOFtay/JB1VaHqRhLu+OaeHI9T9nE1Ld2Y2zO7TtkaBlWL9u19Ro
zOtEp/QbbNws87N5yJQsX15nA/5bkS9w5y+/qCHVeF0QNbWa8pJ7Bg9zLUYFOjHw/knKws6XlPw9
o1TdA9B8lRaIbVrycmCA8B4ywXxzGFgDNyGE9aLGZiEOt6//42L6Ain7TtxVMaHpICN3yfm2O160
2SlnsoQ0se0whR4DmaOXd/13HSU+bQlhy4VB5THWxqXDit8O8sDAZ2gQydag8ahOokaBG0/tr4Hs
9ld6ytBFoiAqTqYcjZuOSea37ipBvdptytoH4GdJhXWILTXnTjGc8bRsBxdG1HeUrmjuPtn+Ksmy
9eD9Gds5F86TW5rESF4Uq2CmO9gtjbzdJRJMWy1XQPRkmwyWWKwS107P6T+kgHDYCg+gIRbPPMQs
X+XYuxlHQ4rj5/BNFEaP6S0MI33Bly0lH2ftOslSPkaYETb/OnoxSKUsHAuCjrT2zNaRb6dOXwST
tZGfsyAKCp1rbTZTnbscBCvL2P/xhhKEUbu1jVSKU2m/km5dEMc973oiM3zD9D6LERJzLpV7yzcE
T8jSJcg0vJEIyKDyCV3YqJGLkewwZLSSHlw/y32rE+baSbALIiaDXrqEehmv11LexZW/6SvIhshc
EC57jaWQUsqOWXQHaLpNtEOBBlDwpyVr0EUmndxk1uo9/g/CNn8ds/8EyShAq4vi86CYmqiGW4aG
zDGA7P0hQBjBS/UOiD1y9/RtsEjGL2Pjs2VRGzGghbTsyHT1rQpjM6a0k2x06rj2v2K9WpoNK1gn
PAqROVUzBwnmVbvo96o4XN+W7tSZbb0Uj4iCAQIg1Q+drO0v3KVkqxEhHkPnL3mL9e9fKP8Yhz5v
qw4/ytcUy0G/Poyy+E6zMknZqguPvFzRvG88sdbI64x7L7I8NAs3USh56VXcfu1pjRNoyoCJyuGM
rQkyFi8nYPb0rrxuqQWAGQESs97IYy/eH6BIX7HPoeHRQUFmmlWmMUo2uuih51R1OMqQZx3i2cQv
+eT5KxUApJQZYTpPj+6r5EFEtM74n81PDVsFJ5AxVMsn2ycFyK+PPEPG7r7Ooju9OwbacUaQW433
PylRZtcKQD3QJuLY5EKw0rb+L2yCCBl8YESXsrwp4isfIEwxS/HuprmRbiNh3owP7RLArMZ+memc
cEcY19bdKHOK3QqCBwDIhc70ShETw2UHrMcpJ8saFNiK4Zmm2+6RGQsd6sdy7cgP6paj2lPfEAR9
2Do1EPkeQizqJVks9aULxiG+B8i+5ILbdfCeto/zqOhxdPDD91HAXwws6S5YBICLUGZ/LMkL6nBm
K97eWfyLX7+tNAFjddckOKgadG6zcnyqtMgiNSal7ZjfpBF8WETUq7NkNL3zPtkL3yd6E4Yz0ZZ8
m+N0KkT/4sgreM2+t9LuIVoaeMrLJGcW/xuZKL5gHMES3h2cHuTDX7edbdBkh12JDhaiQ2VqpI3o
KadS7N2eIMS5W8YBgRTUrRlKfM49O3qmGlJuHESmJGs5p7Ea4jsxntXxF7f8gPeCVZlQ2H53rqg5
WP4dxjDMh8xkD6qlvEBs/bQ38JfvVw6sIJPldnhGqyFcSl9lB3Kest9anw2qpOJoIE6qTp9Pj3Rw
DibMdKsw3+otK+Ky7dRU4BNvnkoitjlUzKohyFkarcMh7MQud3pR8gCaOB7FiYLC8o5Zy0lCD/ZB
U8/w0xaNIoXT7CBtEMqpHGAltfJOI/Qq939nF4Y4v76UYA/niAueWTnpSJecW/Thfw1gy38QolPg
egxjaP0luNOEKbONuXsmOXuLrfTjrRUCTVvhEk+ecz/4mb2XhExIsMd0Jmds+4xLymW/nT2S3svY
NFgig2ZTSd9TXlQnBG5N3EkknIgWk+kLGTK+m1y5n5WhM6ZXM9qmg49ukRuPeL2b0Mg8dFAm+U6O
TF0c6yi9LYCxf3FTG5E3QgVddWiQv7LILmVItjzDvsGDTFVQ3YOgg0ZoA052PG8cG5wWZOsgrUrP
B43fTmQ0/4Jwa6dTBkwyNiYiiepI+9PXq2CNeLhaYJ0VGQQHWIURkKfGipl7HrTT64L9Di7n9VGL
Wrs0LfG4cszCqfIs5cwJBg4SDh5rI8t98YCGzw2VrHKyPr2yPLdlv+ablzGEG2yE3+tdaTa3UpWB
10SfNh7yPwAAqevYadr/mYhw8i8nBF+Doqqmrc0WUSQc7QzZUmDaSzplRICKe2bjoEeXY4SP1qG1
0GhKgfQZCOVlIANk5rzmbHkBHxX/kYuFEalHFIOMt4hkjeBHEwtxcK35oO436qjNQwswwjEXnZuc
H5EB17hqyJbDKdZUfUO5Oi58uRVSuV1CgeAkVcOr0Blt5OpwRnIjkQ1o7Yte0+mNF8/5Sjp5oMkC
NROwJp1NDe4uC5YohIXg8UxkIPYobVzle6+P/hbBFb3r50Y7/QLEnMIiAqbzXTw/JmVoVoigjLFs
Skn+P4WkiN3P5uAzLoMzo/MTs7ge+omp1U26xA8tryTSkGyo1HDMOm944MUe4OFgDu5uiZF+RYwd
eHZ+YFR2Yne2uMmbP1cphk5LCYPtodkjkDVqZh15vOjEYHGvCZXTpB2+eNyu22cGjpHXIRb86MhZ
ncIe0faYLGEcfeyv3nVKcOLYX5HiN3ymqfLtGvJlEgRQnWBVk4drxM23KrC65lBUvic3CXkBK+oJ
C1ziwe9aETqzaDJ7p2TEaK0HuP4LvWVazucV7QUS8/t2EqQnfuYljLCEKS4I9jSJZPjexlQNS8wG
fPYF7kVwawYKs5wX+VDj5sq8oeduP4RwRugSG9doDKaKgSib9l7gFFlpbrjORp8dqAfLNS8qpUsz
8/A6C0FidX3XRacjD4yDRNDkbLcIZIb8MR/K/3yZApbPJSlxoz/KycgTUQj3MB96tzluRPIgyOSh
NWE5YZZd5sDCEv4g8KxADoqQAr02SKDHn+CG5I7mK6OP+PDyzAP0y2Pl+ihvztsRYtd6EdxFy7/q
w7TlS8x4daLZmiAJUSvVJC8UaevBAo4GNkzWcVZxBG6D26ujS712bKrMOKJ70kBdqtoEg7RuOD/U
rFvTmBCdyjl26qbB8whlBbN4hoxdXsuk0k0zTEOUMbEuBTa1199DLAo+IguM950rB8LwmMKzmrRu
q8kcbVA+QhGKobPExSGaj1LHUezYE5du2IfHfSaSHNazVnmD/cGgJfKivAPoOgVGKEL75eRimOVw
7aPD/M1kJJNAaP5UIC6wvtrU6PwcUqvPZE70YIXskklAc8QyJoaZzWM/NLmexEOxvoXw29vadplu
MPd0YtdR4FjgpvNvmZJ91cJKQLpOU5HsqSVkIEfo1CvdobHm8xSTeYfhINC6TFAhobflX7FT9EIB
HfcawPSbHahG5dafi4NfQZRsssVLyZxtVIZHyNIDArDuKKif9Ie1QUx8gZfsvlJCuZyopuW5NCWP
uHujsbxGCKAp59I7eDp6IIhIQTMqJ4q43pTG8HuSvtFCTWafHNkMzfefQoGpHrijkIzzmzRKScqE
HMbHCQYXAjMk7Hg+4J3F8q7Z0AQFPRd7ncrvBhoge93jC1PuCUrYiJgdFETcGSbEWxTRvKXvIB3B
juRa/70ZSqG3P4a9DXEtX8ZnYfUw4Dpc6fJpAUltvnNqivHBe/eaLMIvOT5GpnBH5fbzcu6E49h3
eL7956v0/QX/+B3BPXd8dEAzRSb0h0TkCsYcsAHQR/yjZQ7+eC+/sLUgJBwDKqSOORmq+k2plR0F
7Zrp6at9IyiMUsiswlpfr0ivUcN2wZCAxAZc0mQO9OLauiiC/BLa/SsZSm5RUSnhI1JqwWbMU7j0
yaxqsjhzGtJ6bJrJXEk4DBhdHLPmKh1ht6jLyWdCiaIkCNahJM9fh0zKVMhkr3sROaCqg/UQgpSU
aNHDw6sME/ZoSFE2jmJWa0cw4amtWP1w8ONyUXut0HJoDlKRP9BpSQBqkGfvcU59g7ij1EC/xQ3P
l11XvMVBPS8W36sVbKv5V2+DotZEV2cxigSTyHNZ2R8SAcWhLA055EDGXfw8D+vPsxRnLGuqAaVU
ujjX/rx84Qd1QwnUVoVgkqO5ZN5/rmPK4AopvUZ6k2XvWrTLl5eknjYIrBr6ATWiZ39+JklwCOpS
JpmG1yVdLWyBl4ghenstVT+VdZRw0bZJ25zkGV3i14Hw8GDJ1/2Vu4VBfjguwXoLWX56GY45LrwW
sKttZm+BTHYXskTTHu5QoZ7vfaxkU12kv3FL35vMHCak0jyZzG2BbOlLu+RjOjKKmFugf0LjQYCg
FSE8DhPp1eR7FlKjXYZlJJ8mjl0hC53s2VWd2QJoSeO/N7Vtv+Q1H7AfuIe3YCug18pVNGBoxaU7
BcTAHxVCZhqnROuzLPHYgTMoHpeQci5eWrrPT8Dd7RDLrkRo2u2/QNq15TnoIqx0LdjphMd3rf6x
mUAkM8Geub2DLSST/W0TJI9k9EAWpUODuLQ3DpPN6BXpI9pOuWV107VSqA6YmzsVU/+syUliMDfl
Lu43+PXE7TBhN0IgoTtFJl11ta7aZeTVLYveBIXSVhc3snHFb369GqZrNf8f5kDLV846wSmTNwO/
gHWTLLb6eKLNWQn90gYjJlmyydK8GDPMk7uixMfBPQI07s3bVl1ingSwFDto2CYcFZv/tUJOlpdr
udOTq4Zn2oO8i9iYD3DLh3ctAX1dbDw/g7PwhmLcbmflgkGHGwRoUQOWr9tNykLpcOfAHj0P10uy
wBQLQx6iQh97IhVA3uSN4dk4Ota4r+0bXIDnD+Vx0/B21StV5xqT0njC2iyqm9gPChukkLU7YdVL
67uyUIM18p/mVMCw6Tg02M4xUf6j8S+sgqiowR2nnQprHnxqSEu8nKFyyhurL8sf20JtzKZY5Tav
tsvzqixpGDM4a+LhhicLv/3pifFGa2uhOvhVNCEMv5OmbBBYwKsjBwLYyxHpjx1z6d/KhIm/u0ZV
x0/aypY5jJovdWFqMEJ8fqeM5/DW4zX2SY8NRBWYZCDuiFIgz70EKKfTcW3iFK49n4AIEZcZlz8g
SGDsz6TFKP9jtre3VRnsOfWpY0zJFP1nEjLabJ9B2C1J1NGDCClwHDG6Yyhx6M4DTIk5cotsdM7G
MYmabqbyehMqojGLgn4Beng0NYAdwpotoXk9ANoq0CGVk3VCEkVJmIoilrPlHLhjq/OTmiwE8u2o
1QrIBbQ4xQ0R53HZKc0GVpE6DRiI20JGwLRkiH7v4pcaAjL5ak3G5etP+rZ4SEyGpvsUVzgFNBdF
jTf8JosbPxgRb88PSdZmg4DixPajQGehxQ/IH8SJUtkzvHBbZKGDZGYXvnGE+brW0+fLMNCj/YT4
9bjgqggPQOStmcrGqXozooY5tyeJGLZdUUH/1b95AOhD2GpyJZgUnbOhaVzqcee6VSjRncD5cuhb
IM2q0hfsz+iqyad/GYmpTTZY/MJeFz9jl/b22QYyWilUZFesDCb6jV2ermlAaLYtDw49CI1ZaAxj
TGvwhSyh3uF2udj9C7XtSAmN1P+1cd+DEitB1/SF69PNNHSDhq4BQdQGguiHRd9BwDRVln1dH/oo
1oE0GHJt0JePGMooKKgxrOtC0crF/AYXHu5yDFuCnkI88ta3ZgPBBGrcVcid03fbO1EUpJ8DxyTy
Zlwiq5gNPCCzp2/1S3ov2x4PL86BFdaoCBfPP8kMv5yW1LfoWluO7ota2Ip9rCp16iDPw9WKMIa/
h+HO3x8lJsvfwpmdc7d0WFEv1EiMUJdWVi0Xh2WheEZhbJO3WrNRYNlQWCDI5HS95Dd+d8rAabml
L+KwX0bkoptV5eEpWz+HkEbSDSBUKAjWg9uaOJnc4mH+4A7vNSOOSyG2XN2+zp6P3rQlUvrad6RW
usOPGIw9KacBoq2RF8z4gb8reuaHIo5fA4Tb44EMweDRwblaSXpwjQ5dz8XH8tCftyy8ZkGBYmVr
Ccvp7B899I43ZKe0/TR0ox4AZ9Kw+9F4c7aW+kCihF2FRhW/POccUz0Du/wrrw7cESWgfYM+lySP
cWRC4FatKGn7v71W40O6SwJwxWVe7hiiczhVPcUKOHcSmysZgYd1Z2893Cjiett4O/3F5OfHSNEq
dCE8HczQDsXITqbKYYq+eIrSHGkhXTg/CHRXLWbFpp7XH1yBuLcdU1tti4+oIpzBGZ0kYWDS2Zxj
+YOaf9bQJTefQb37DXzdFaiLQKOvYpqdbCjI7u+0KcEucFYpyRQgd6E/l7v5JXkcxxNBe4BD3r2K
m1C4CKC9cGiDA+AXEAwToMUusJzA1PC4xMDRGeJcSdDrW/KnX+B7ATQb7nrRmV7LgoBNZyOCuLEA
8TslRr63W0HaY/pq/L5IDbkS8/ijZcyfR3cuo0q9puCtUwKmr4XHgLtq9i86AOxrXYJbiB4GWUKu
lAZSUXB5fG6slKuhO1SNk+eRHC4zOLRcKFIfQfE6a1GFdKgBlntoBEy6z06C6gz8OiCFV7pSJrdW
U3bFWSyHyWRItyn+cmRrxwFMxUm8ic2gv5h6e+6joL7+zNuvHGCj0C/to/BqLKNxwfP03a3n4sTd
MdZLO7bSrgegAB7GWAeGI5kykpclQx9bozUU5Ra2LO2Lhn3BsUdyUaTWyFWkTS2HTQEowWVVE76b
aHaS27xOxN9lgUnCcNOzygeq4cuhI17p+MsiUm753igoMywN0DLhdMkFWCYWRAmrUyCjl+Nlh6eg
qIChrWv9q6U7Aj0rQAmTW3s9zjotCNPYN4tHchxBRTvZ54HGPyJ0bL7qwls55hVKS5iroWtjMDDN
UrKBUuaWMqx3slY++gWL/k8vkOghIQzUS8RiHpF0Js/oqNTp6yJ/GTtoQ47r673usWyoAW5iRxAf
2vxOF/3lX4EC/Ljb7h0RxQ8bzApr5GigNqQJmdQSdZvwJ+OcSpNTdT3EwRx1W9gCaLkgRWZP1zsa
vk7+LYkF2n0aIJHbIAJc7AnnVYp3aT0L/YFmVRzQ25FUZ3VeWzoqZH5mJiPFLy0HKnhUpg0nYPV3
nK0naCQTmyXs4jyrQn12EA5G7/+xGEdDiu2kUG5OFTvwKopEpstORQ5bgi0VtVQs1PCbIeqAFWFS
5MiNs6Sf5V8F5LBJfqMhPmpvPj7oq8yJW7SKDYheg/LxyitG2ck+8+37/6Fhn4KldKrRKPc+ufH1
TMNvkX1kHh8wljogKL2oCZQ1rAFq2O2BTzOEbInBM28/PqqqgzzUOP6Il5BugpXIUfvdSUddRQHq
zqv3CdPmQ7sWYckDJmP6Us35KSy1z7qIQLlnO/76ntoVpxy5cm1sOrziRX/mGMwfnf7Qh71rdAo9
iMzfCYDdv5I8/CWEddQuMICKsRRO6qt+tTu2yIpUh9djQP3SzK/29+2HZOMMSW3VESnDjFZVoMeZ
XxrBpWQqLdMSXZQpIcuqxvfGreKmBT892TrE2JrmzrSQ5IFp/p5v3jkV0gU16XR9hgV9DTAi7+OD
IvAhWV+f+1/cUnaPhiVD5p9Q8/Q8fSWp+Sc8OHDZWwp07IMvMP4lPXEgXbSgT0b6wX1b5ofjREgj
Gpz+HfHE/y6YLJbeMTt3C5XPHwI+/QgB6y4NfF9nD9+qX5RLfhHxUgQsEUAwH/W7VLQ9eWgOaDcZ
UYxhcnuynIIpXK/8Nh/7upr+Lt2+ZQ9MXKqbya+nph/0Txn4vTIXWryx5/vnusk4qQvCvpOIxfuU
szb64PfT8rY+8dgFs1o0n/jgQrGGrXjM5RV+LwFMFQGU8EJsb/itwJB1rvECZtV9r5Qfpl8dG0D9
z77+1y51pY+DAmt/15zLhOMk03JED8DsYdU/20XVLr4j90GRhrR5EUF3BX8SkijCgZfZ8jF09Uhs
KQDi/jZHSYi7awMmrPFwSO9yJ3Ammx0jIM+D33CAUpmT8ZyoYA5LQ63nuDwbh52qqaYLmDGWTXqi
wbAd0a6YgUm9tLUEEcO08X+nkTfwJWhq3Vy7BTuf4XvGcojEBV32eAVcAC2u6jyWBz8OoGnNU9NF
4benzgJYk6IaQ0/CgN5ltRlg+dacCTeEFynTLOL0uMLpIZSNAmmbYEd5Aq51XUMZdBoAuNRnK5rj
SPFaq5XZY3MJ4tED472HukOJaiMaOtfLk71YXWMqfYXI0R66DpZKvHUdZviKX//kEex4ZfeloFQA
IDkgT8hZYPsJzLVMf/z3J2ZgZkUnHd1gEqcoe4SVkzpoH4Sn1Viv4XjGnWBJ3d9NV+aYgMjkaSyg
hgggDU3+fKutqcjRu+dsg8L+CFrnwQADP41QSq0x6m6fe8cUTLH5gl0UAEc9R26Zhe2MkY2Lu3zf
TaXZeX73H8oDTcfx7jNRBXb7oroBU4e1cf1hhdvC6OBAPf1W27xKoddnxT8tjXUq/FlChe0iMeRE
O93CmU+n3kcJzvkpc+gHZhaxO6mh7GTpGOZuxXpBUI8XF69K+wFEng9YQUqao3z/knDwumpWk3X+
FoRDdHY8my9NnUWO1pZkLbj01Ew+SxsPvohvTFOQBtzrqE2Qm7ctkYfvgRoJLwMkcXkzJXv54mGc
alx0u25Ee1cbqXzGasozFhWtA+yLaD/Dy7ejWe5UrI144/gcf/A9gvGB9gq8xD3ICOpIXrLvvtRj
Bdg6NjdqDiExJOy/tho/cilXMwuEm5cn8c+Fcf5vIzKNrm/uCnAaWmjmJpsxcO5G61btBY1KkkYh
D/XW14NqDXp/gP2p8l4g3YZOVDYYi2qA5i46A0psDNVuqoNREOZw8G56B+SvWkC54NpAXrI+Sa67
p7QqNhndy3sbFE1iRTXy99liOFEvb6NPiFd+sutS9olxXWdv0e+Dh+WDUPnCO+T9Cu9xTg3g/Rid
hj2feMRKtDDxxYMHwUfWosxI06/+R3il161spHGX34lJ/pl//Ln5OfplL9q4Ljf7RCDC3PHD3Z6x
vI0EJDWmgAdRJrgMlgKylfEXC8IQcC51cjpmH8DTpeKBarjJjJiz423NwfWvTT7sBapw4sg3JRvo
fG2iYoydrhunOFOLAyYIGBsiFfIEWL4cKKuhLohEjvHmyBACNL9/q2kaCJ3XNpEBnGkNeREE6jZ0
2KRD1kp6xeO6KDfNtH/jsG3mFjyf7o7nfzu0XRkA6C7xNkcNaCbaHBuPCFLWiu7eAUp/Ebbv1goP
wPqPrtcdbfk0MY7+K2ZCau7IbCxSroT7c8ZuJZf9Ui+QorJWTBiaBuT7T3InDS6PU1bTFBt1Anq3
r642z97KyA5TLVWO0BrL5RnyRHcpW+Bav2ZHxszNQe40+WVW5KmsWV9SMmwsAZ/svrXflzz3SoTk
CvMetrAGPotheLrtIQ5p90GNtMgWfkhHkLF3qaRPzjzlisS2DmhQF+cA6+GXwrd7emYfsB0TXDHo
ThUvFvdKk59bPu37ipYIk2THkqIRhHiNqELmBfbgoU/FBCGOSPn6fyEB4uw/gZhc9r9s3fv+o/gG
DNp/ZYlQ0j2yzkl7cgO0hD5axdnXqzkn6OlfoXhUjn8pYv4qu+uZtNwTlWo/rRDtETuWb17yekf3
KA5RCu8oEQqdT6G4pIS6Wepsk39X7x7dpHT5+EjPfbHQzxMeO4M7l/CDkBV2wczgIt6JDKUhvOfu
UMBsBMMK8wYx55NdQXRtgRziWGEJRMXFOAVZRLm3ICIvdQU7oiTG6/wcM+M43M7D4JZzi6rcF95o
tgFIG/sqRqQsAcVw24KceSstqPO1Yq4SHahGN3G4olIJKk+0cG8WPcW3dfvKASvQYJyTyAn3pVDW
u7z3x3fS+7TKC1RUcHS3h15d/9QlUqu7p30vcwnHwDFEVEMKRi6vP1PD+NmcHKaiS5bEpOZmLVxE
cXomP2AZEMzo23Bqr1SomN1hfrv1kliFad66+yrHdFaHG+cRlaMaKEXrgKPWkcQ4q0PmSg9Kkx5M
HPiHxgLLdl5VU2fdxWC7VpP7f6Sn/AKmt92Hk4lJyYLlxTi2BBqBt5RURFBnfufPEo7c+EDZUOw4
pxlvbg9o2N7vWSlgs3qVjNuMhNW59NCrXzgf3gPbrocF6HTgPbjlUxemz2U2+V9dB0JAF7fyU9Oq
itP+nEbM0wZZAtNTHDsI4sWBv1vnitOKqbeaGsZ+0aBX2lVS8dld53E19k4dkLiFO8RAMDkcV1yN
36IXmY9WkFf3V2VgKdisqTzG233AVhoGUDSedIyO5JL2v3wt7pbay/gr1J9/st7W4FcjEX8i7ZcB
PrbG7DEv0Z718MCdEYvz1U+1fc6oAweAzWYUqPcODE8yviggtxVBVpGbODVbykfnw6sNCwwdSteV
KNSEPBhfi7qp90oGyZS1t9JDekC2EDJc5njqSjCYeUqjVwE7vORHUSR3NUy/KDPaX9FUsmsJbrto
iqirAuG3EycRMVrZ9w+kTiHi5+/G43wMa9QuFzQ1GgZf5AF75FmadK/HaS9fs71wriCdBwaPGz3J
5yCqpUTrJcy6apqVvLMlI9gA3y5Oijw+Gb7DdJkDLsQGple6k1GolA1qzlzCMzDXbHy/nXZWNEXs
VQltdWCA6KUH9QCrhPGke7htKi5Usbz2mltNRP6CIqS5J4mVUMxSnEDP3v9AnopHPot4b/QUZuwf
meX1vLnZKH/yZEK59uSFrWmrEpxsN5CIK24JJ3q0axK+j65tH3IdYWSoKe1SOdGZ/zKbZfvCQtek
NkZ3BsFSV2jFls8f+BRcg0G0srBvDsNyeJBhV4TkcJcn0dLJrCa3XoTit4BmmSTvvm8+D6/1IX/f
usNkmByUFwLWkr6y1uxEP9um63fR7hWodx3WY8oWyJ5ykMi+BUgVBNBU5qZdVfovNOlyfHfbDJFj
r7R7ssGn5Y1qgqkorcmEmTdoeASwO+fkHs/kdCmNXTk1hKWzYt3qi47rqGrnodOZiBAsCgvlUUgr
TGYSbvKlltFZ+0p3kKHOy3nBwLNB7vLLpPXK+wK2drDX2tVnv7tTkGfnEf5jLGuXWVCkeyeoRrvV
Q4k/GU4ijbg7fxhC1Bot3OovhkCRMvCGqbub0nte0krHAjgfkgpKmZ4Wa4KE3EDVW3RZE2rNDwv0
cbK5Ys6fOIbBBtfZ5ronRauoeiLuQVhv/H6okOaZMqAXc2JTXAiV8CvbuYPr0Whfi0yQOYWfi+fo
XQEn6nPvaupwbOoUltpgAuEH3z6qHLo0rAPh/E1f4p5lN7SjaIBvWkd4+8ksALFoE+gv7TtDgHCA
LnA7RkwxKWn7sGUfmBVYdI1S8fe7sDwUGsWb1FR2BsY2GpuTk+qhpImY3AkRoU3Gl+44FxFIwmQM
Q7qBJ7TFgk9fYaPPDg8u6C6Edr324v+G1tLrAFQbKXlZPjxyMrmt4a1goXSVZrmoLnFBz0dORPFl
EVUJeDvKSpJ7xc+eDRH/WYbI/jo5HJXzpOzmIwIYVoay4X4Mm45ZNAQHnv7wvsGbHWSaa6TDMNiI
vK4o5/YD3O+C7kUGqikEuPtj+ZGzOTJzvqgkTxZv78WbPezD7PB7em7Xq4+e0vAEPpLBou5QlxS8
exSosnJtx6kEAZ9QG3wIfneLsWqoMmf5MPtQA+e3svPhafD8sHw1xfpbNMI2ArI/8E49PlTvPe5G
uxQBS3+dVFNfeFPQYHdLYORy0oPPrxKwNsmHPs56YGnVmYOzSP5vYqqBkV79jDGH03XlP3xnP3FT
HpaojqxWwUkzFa3o2Kxh0TE555HX7qfhjigSEAXErDI3UGpzYycLyR00qtZf5h4gSEUyN7YeQSXG
Gvzy69dBS64sjMixn+fv254G4EJM5SNKaZOeFxu9vUEbIa6pyZHd7Dn7WW9zZRak+Vn/UxCdg2EF
DwbCzumUUc15hK39vvcMJydgfV18Y8aQHV5dUdyDc6krIV6Wv4gkKi06Rv+BpS8I4yz4om1oDyr3
zm578Ep0h+D0fHHRxq5gMJRePYbROeaCpgO53oiBs6YjTDlFEIKQKDNtLNLG2pkDCpr2sOsW3x1/
PEj8Pn1hCjyOyguVHKOG2BG6/h8jB1ZZLVBt4w47TMlF6yZvcD+bGiVgIrODS8pM2nA8bLMdO/wZ
CI7gjZh9ObVwf4POENDK4B1/X0EXe7eutsjj5d5IaXI14nY377oZ7jcES/wg1fQwpZw17hnWdSPc
FuPZYlPB9MjWvupDBA/Q/xbjqu+bxzvJA6eQYD9SE+khi4+7DtVxWuuGnWNlJ5cJGI+Slk+o+4AZ
QhC3F5HIOr+0GEUw0POrQ2pQT8PjmOuIm556TEElqyekVjcp1lOslLNst3qFq/uBKmaswx15jT45
JYJFkUU0O4cy1ZtXIijxNqGbDHU/sWiLOoht8HJaozNYnYE7WKOcj/7YZLHS2Oladk/72HF83fyi
pzW4HxDNQ5gWj0z+H1dbW/LwUlhTx1MwBag9/65ffSpQIFKN7GCAzQAG4+LFJpaJ5G1giGOys4FM
+0kRRysJmXbGFaEZJlCGYiGd1AAPbkSJuChOU0/t6rk/5ttozKAHgsPArwxGfTY1gm38gjolJ4P7
wbCtNY1IQkYf+uEPs4yxzhPwb+ktUB/6wQ4QBv4FfHrQNO2PuUcfWQy45kXTEW9pCMCH3Zqv05F+
itS/SqbxJ34xTqs3PiJ/dk8S2Mox9CqQPzIfqj0KHBmrU3LTonpy0U6PgHgbF53mJ7+RmbefiLT3
pvwwKsanKh7cyN3HnNtRjcsDumE2GQW+OG1yJZl5VZUi+LSH9rzo3RPbPwptsUXUUfrLbJMvBNrg
LrHUrXNP+zPGBxJMfxQso+Ba2vcOqmmvuLycKsB6TZCOxDOwti/ssmNvGf8XI0KVJZYr/bVpawVI
Ui7AO8EGWHFxKn6at8eWTbVXgurC3bTeTUu4LYeyLAQCWt06DgdcALZA/5/TKKW1vWIu7Rp0U8LS
eQM9vGLQrJro/xKltZB5vSrOCKA5C1OCu9TVkVUuY9Vnp+HCbU3AS/qUd/hdP9kOwjnn3I3FFNYL
nCy/9fGxRncHSdq5J/7vHlYrEmbD2w15nVhw0cGnxreYf/TNWDveA1M6ieDa/lQ5TGF+S3LO0oPh
35UL5CWG/Sn++3IE0GLcFgcCamDgCLb/LGjLzKRdscnqyRiOOdO15OI8j46E1Y+eNi1sZ60ShisQ
4EoG7RNiR1+HNBK+y4PsW/43lwuZ3g0yhfcIeGL1BpL0T89EiCTZcbtDcFUwbNHpVCO31a/ObFcC
DiMNlENgVAHGUlDwFNJan3xHsND8BG5/yvZmz5rS2OHRHRDOS2ud15QtS2CUP8xIWpVGwY0E1btN
jN/0iCb8yxHxZA+j+zOJOX167OgaIFl64J9n6ESA2cDiokHXg9uebQsLr66keFUd4vEdI82fF2Bn
FGtSxTQgiq8R/3blTRuGRa1nEmZyKOnCSkVcYTzUriGkrZwws4TwTC7CbW6kk9FWlvL+LJscBw+s
/Cuehrz3okUz6sZgPSoxEj6WvspEQUxx1RNR9xIJ9gcqE8n3JwS6w/4SEMAwvgvXbGw/sWUQVj72
aDEG28BsU8A8cNCcXTFQx563b0ylxj2KOrC+EQWo48NDrFac+fex8rGmToO7cJO6d36u3wFP42DP
yojp5/lctezzVtJSjavnwsaouRgCe+yDO1/JGpVeRvox/qvH/UrXHl9xBe+L02QgSCLuWx8g14qW
AvrDJSgUHK36RhznWlyoQbs/TG8inUwp7XwjJ3cBlXx4qKtaXO5dvg5TKC0q8gXkW8UeuCzM0wNT
9VKnkbkJeeFztbIFVyK92ZgoCWfIEYOJuvXLuwXRXcP8rDNuOhZFPLS+qMTkL3zLX3AKnULOZtBQ
+MDTujmpvdhK6TPcj1WaY9GvQtnYTWMJrvtSbPpZkADNnkb8nPV5BLI+v2CT1PfAmGo1AcR4t21U
QwP8Vcsy/2+j6f6RQQC2HN13qljTlcP9Lko/JzzB/tGgnm+WyXqH1w5kOxJsb9XlOpYbTuMnGhos
MJ/Enn27IDAU2W5RVv6YyoVuiBWZ8BdZUX29FlYyQDB//JWO53+zicPcFdDNjjGSAc88p8sMP+UE
SUWzS5qOK/t9Ppk2X6SGxXjcL/HqxdU3KMkY1z0QH734ZYfSgeOGbkSATfwQwWC/slGMwCv65zCh
ZNw5lXtE6DiqBrfrsLdmYjrUMxPNVivm0XWx5uW6CZbq6xEFX16vEFtChBth992C/r01GifPa5nf
zj7Q6ZbGlVLpEsSskRqVESKHhqVcjCr1MjqCvakC8RFdA8VydBHB73ZsXL+ob+Y7FgB7mB4VHe+9
FQVzO8i4D2ht1944uMi/LO4REvNH0BIxj7diNLCxBAKLVuQaQsZzABaDf3nACXLBdnJaIHtoK1YB
n6p8L6skzTqqtISqjkUSq5LojkBwADiMBi7i0JVhbMGk9QpSt1crSYeoPx9WQY3gGeShpDHAsYJs
qVjYOEGc4vuMj2jz4ClAk84hW39QdpSG1Z2PuQidP6sqPKAtbcBw8EAU6Jg/LoBSKiSj1k8IYSYF
+Nmi6GkvKB3eKaf/oyBO6QWVapuuxRSZ/iNB9+t92fkx7tw1udX3HNhLtkMhp9ZAz9JKzF0N28Sl
M6PwRFL0jl/+BrJSZGqcEcUzrLqN5NY5EENeoARit2aUGWrYfbqxma69ZoJEO5LTCkC+QQw1p9g5
/dfx9J99PiLHhexG43FvAL2qufgAuPsUU5fTsB/LpKar/U96k2sHO9V9RwVBTdZ/jexhB8+BbYBK
M04nrMT2zU11WPKWEUlC3gOXjjt8FAmEJgfKwMqONqAYpOBdGTiYQfd6ru2+YhBZ6QbZQiNtExER
tl8zsbjv4UkpxPBJKq+7wBEVVcM4lVj5efT7D12QJNguLegYMxD/hKSkTKgNt8aNiTn3M7P/bJ96
mV8AQexyHz1GzjYcesCzjGC1gNhJ3CKHLED/Vpqi7bHKK4LhEOLVre/YBfM5qXE9ws06IAvWZgLg
nkHS1gjzJSo4++46FMi8ePOCMVBy3f47lpTj6f4+ba8MPCsE18MYCSKZUfXUSlVVH66JUVd/3/ph
jpGmh349wvf419shnBPgQdsPRk7oPZDXm+8zk8IK9XDpsrbWeCdyavcXZLoe2GZ9wZP7Ecr0i/uP
OtefGQ6WjeKchCQALEy4bxr7hrPh95cfLDK9tzYXpLKfd2GhmKERq/DBd/Kpplmr6Uvx6PR52GCH
PnzGvdGN35roFFE7LZSmfKuult3rW03x798LJ7iv7cAkosg6VnI5oSv31/0txIObzhtuAfi1qs4A
GSMz75iJG3a+Gvj5s+2GzY0qyMxC+ouy0Fy7eD5ZYlCVLVLBMtJHwXZsWqrllDhx59zCxuyYNDbC
h3ZELGubPULpj1bz4NDQKkvwJYfJLiwkbcaaLuIc+k6Is+dF7NXcx4SkGR3xsSkv1htwUcsvFM1u
6ukizrMqYrGEEIoI3w+Kntn7ovMLcf4YPxB8oRWRBzSeKaVjmov83yNX1LuQeMPCVF2FBh7W9k76
1ibveGGpkQQuH++52yfS6BzXpL8N/yp0koYTcc0ZvMkmJW6vRk+qiZZnCAegZnRKf7A5+jPp+mtp
x4zUPPZwb/Knk4ETSLOLf4Tz8Uy2K9hkHOmgzB58dO/Za9jmw6QQtjNxwPYSs0aFf2nn6du7U8p2
HT+HUvUufdf3JlMDKFg1zgHsjSFJo30qhPjZ0Grb3SPB8DKjsFS4n8KkhOOcxYwFyjBOd/9F9rJJ
0gFsw52rlCpd1HK6BtAsQu5IDHneV8j0+uIeJIDSzjuJ1G6E+g3KeHP9IXABs4b+E2VwRkVTBPSQ
+8O5BBO/1u9EdrF3aGRjuYRS3Wq6yg7XoxyRKHm/ooMhSTBAr46JducVAW44nq29rWwQoOy4uzFn
lvt6ul1fP6FcM3Wjl8z6UQNyIasxoWt2QpVfIM7z3XpmNiZBvP7GICSDCTXUbQpV40vq1rV+3qhe
YhNHl0f4fXB006/wLJqHwW6HKINqi13M9O27cCly6q4LN9oor0CFzZp5e92IioUQR8SOmOK/c8TL
0KNSH5LP9Rfbu0WlZDqAcQamrnu6ApBjKFlwM3TDCs/W73Pzjy+6O/BsCBINotaw2VXcf+RrWzFv
xyeBLNGVXZ5OeRYG4Am+uD/e3IzxVVMJIQAzdLPpiNMBuX/j7qwCCjeMm9rMZsEYJgIcAUxw9J/N
E7KVGlJRRCNW+nbh4xvmBHtidavcsPmhsll9aZxyMKQCh4geh8fiX9FeNElRU7OlHcih2vw3BQrN
RwthZ+xp3SrqMsuebku1F+lq3PFBWAeUwf2tXfLNz459nfeMWLeptjdlvD6sAXe1Kxt/5E7CdKym
U5qEd69JIrpkLYgfS5TMNrqcTL+/bECED419b2czbsB5lZ5pYecJ609NPhirEawFzGjAUjWijrEH
TuAO7Q+y/RC7UQb+7zFqzqNuCmu75WBsOd83JTbHR7Dx9ZnIP5fRWjYj6JqqICoGOK/c7YmPMXZr
NW0SO44LA52C3hBG5/XGYCF0I35bCVp6r75rMVOA0Eq+t5iEVOsW16+r1+GjOPRwd8S5vcfgRIkb
etNMYW9j3lwIDb2VPXxmtfgzZg1V8aTb38UwHQYgABcktamr97C7ifeo4EPoa85XViFdPHblta4t
sSlUJ6HilAwLT3iJP31pCcg4He1WvH9lHt6m3vFxYaqsSeADXkZAPJRy6Sn/o7mpLY7NcvMqmQAw
oqVvdvg++1e0uU4yhCh3sBqlQ77LTRUiUCncHY9+OOcEiU6Jsf7xgPaztCoGWbATsh4YtBAfFmF5
VJz2I8UkDXMQiu9yxh13pFqIacauIM7s/UsVOPtJd5z4l3cvovL/QteFEf2IHEkolNINC/XY3/oq
iutgn+hmAZpNGybDqoVIa9c3oykC+E597zHmaJkE1FKSu082cMIwAdP01rfTJmChRTGWfaDMJhNS
neahKdDbDM2QdB0hYc1y3/d02ENP4rRqhxksu73Tl1Pi75SM+OvNlJvzx4fN1/Tcu2E3NoEoLX3i
2eNgbAEEAgVzpmmDkaYtlJAvt9rdyYO4uVruPh75KyqQRv+YATe2jCja49iFX4aIR1xxn4EnixNw
tR+FPQCRJ+6335ug6bvJWxkuRD3/rUKo3ERhDn05Ctuew0xq9wPFqEZmP78x185jpq++E0y2/lhL
4+XkqobxRmDfPLohuCKKA63qI0WxTZQcI5+6xjABV77AhYa59mQ2hXb1Sqb7xVhu7+fZ/mZh+/SS
9mf4Ampb4rBoD6ooPZXaUKK7RaIINj37HV9fvkJtxR2o3eOMV+iEXDyHoc681hSOooORuN4hGGmM
MQevOHaycDj830leQaH00476ZM+vaib+ytCTtEMt2FjUfkU7Ap1AzXUmTEi1QG9jE1qAhr7BMclX
UyOmbTLoT6jzBDWy/YSqbQ5L8X7Trunip9b6qKRj35Ga9HdBJ+GE8ed+xKtk4LTLfyInOZJ+QQ+j
sJcCqqZ8UVG/JFXSoLyUJLD/ee82xdLr4CkAeGDRs43hh7lG83aEP4wtorLeLBtscYsjTvgNNJ2A
w6xwP78JHuegcimdbe4iMd2OioKYyyCPLCfIbKf46R1PpQgyLtL/cHbWkvK6p4OQlAbsmJAP8BGQ
7P2TDhfTm2S1o66V4oD5IJfdR3dCVbYJNmpjTbKTqAI0m1kRxa4h+G4/YVD7ctWIDW/65cpuo5cJ
BBg0avFehPkpSPIId49kIHiOvZKvpfegrm/xJhbEYc1zCyr4V1sC6O2mHe//bJi32QhMcy5uW5vy
dJKBYwH9Z/c/DkjgNhyWaUN17WAz8BIrH7/KxldGntjBZvvwA5i/IE7reMJrHobztLMoWAkjgvGp
EAMKJqXa3ebYC1OyDx5YlauWLmzqvGsAss2Q9giRoRx2/xzbBZr4kz7z46hJtE29xAiG1ZducDvs
I9Xoh2pORp8+wf0HUCA56VJq9tjNWfKwkTO4S65mRldbww5hIx85tJ4QCbNSV1XLu+BvDA8q83hy
lwAtXvf9/V6HfO54SVF9eC3irHdRzZ7EAtIbvwq4dOpygs5L20aSaQ1SUWlXSucoQbXAvjZXM5DQ
0vxYSfaCcHRc4K0gba5983R3etdGcqX4V/fdwR56SdRxy81dsVWSiakVx0+YjsZ5leTpZaRUbVsF
Xw3F1pWF+7zfO5u+Pw+pTJWgDmi9f0K57bYaOyv821n8c7EoYAIfRh90ChFmiUcBxviok69GsttB
jKubaMhGCk5KS+/SIKWLNcGHclWiU+wNY0w0t6VF2GObCzRla3T3hfSx9Q9hAPWtzpxux/RJSBM9
4UHVNQ1XeEj6TZou27vtdGgYNhjm1u+G7nxjftnW6Rum7BlVMfBvTBbnFBIDFg0grFoy8HD+WOkn
HFCdxkwmyxEh7uzdD8KX/wX6JXW7I+S/I1Y/nlE6ocya1yFDpfKGSxz7nHq8ZHpxPikTRpC0R+CR
RaGhF1pVnGyp9yS/WnIBTyKaU5XngbNo50YTEoJhyJPoidDPK6044DwQf8MTbQmLa52AGtVIm81p
plzoSBi8lMoTXqpMQM4ZjweNmdyq09pRQ6017XVN/Fe7TuTZjDZQhW6DGCa4ZkAYmPG6UKLc2ATn
/8FiRQjRSa7UbaPV30BpptntkGE4GaUsDcvEmataaDcHNRIPQO/KxvtWE7tzlu1PNp89dMcw6I05
5bgpFoztfPUnUOlJERqkeqoatGvIeaRRG5IaG4mHiX7ilvTWTRgcR8gAC1EKBusGMLneMpM2vl9U
GIAC0RZPtIOLbILq1StBPDj954ku8OUvNW9uKg0UEfWt6tYDK1kA6Nz4CQWA4TOjTReJh4yZv2af
pWytoapZvBR1NN2Djo9m/2V77v/WGRdqSFfVUNX95+o2sSZqMf5j4v34STe0S/AymwLq+dzf/RVq
sSBSGZ5tgm2vo6qrnXjzNuP5Bdj9IQ0gRCKyWfNfR4d2v/K549VefYpIvDYeWnQyEJjZia/HsVP7
F25sz2NXzDKbFvWa12nhDaM7LDBH53dZy3LnHqyqqezsBn+8DhQVIaRvbEmrySVy0ItrrEx5u7Hb
EG4NNT0d6laT/N2H0OjhoNsVSojJEmFp/294iZu3KeuLHXhaGr/Tja2j/bJXcKIYB2M7O2eS0yNJ
PEdaBI70xJuGfoxlWKCtw/ICW6SDWqT22cos3CJRJbxkmFuEty6/ZsbZUX07fUKBZeUCMyprc+AT
6PPMbAGg01o4RjpcFo1zgRO1eqPj2l/fR6dlLXm69/gARxX4a7h/bO4KlRCi3W9Zn8P7W6FFT5sJ
8C39ja82fXBzoctMUhrDrT3yBQPP3qLJPEQ8sDukG0mNSyQQCErzHm31qstRlSLnQVs3LstAZ8RK
W9qZrRHf/4vOtq86CNXaIzIKkuvE3hnYzXAVd0G1mp0PjxFoBwyLlQPF2nPBXqltDqqD8k56yBBE
p9gGaKyqcGNhPzk5dboUvnmNEHrkVIA0XeaTBK2ZulQmQ3h8wguJJHnh0oDJkPVldxmdvxBSljD6
GCBFJ1+4EZvcpiR6o7VAi5VuideE1bU5ewhjOJv0S4a1Db/2lksySwt1R2SYqXJW9LN5xCvE0oZ2
dKCKzpf5VaPKbD08uKL/gu0gINgqKMvx4VqyONLWw0vInz+q4N0s8ocyURXDCsGPBYDbol728RmC
5lqMrE/mI6LNE5iqZZnQVXCptIHSWR9jSl2SrLEgbpZ9KNkHkAXwechM9id9cjizqyFtCrDoTUhV
G9LiNLfEfunEDwH45h8km5o3OK6m4hoL415IeqdBfScKnJDTDSvjDXSjdxuI7/eXPWxQIpVGfPYK
3KiqK12RKN8Qx0kbOYhT08DjEF13VCtdYYmdK/OCbxlyXKgapaxL8VoxO/PfKV8h0dh4aMqlJY1K
gOQc+VcW3+Ro58lm/PYEX4h6QiU3GfhN9yYlagqCCm0mVl3r/r+lQov9l25tmqZIH2GZXB6HJl2s
ki+NnYrkZ7jVZq9rddiE5lneci96hXwuzrtk70hA0wfVIEsu36kBl7E60BwNpsMKy9VODVethuJx
1ktQMxFUp4gdExAI+PJ10YeBOZ83ZcecWC4uZQ3C4v6ocZnbE6brxJQwWwY5qzytMPj5SbG99XQi
di8T5bs6jdLfl1+u/zPSvJrWhuCIqiwYNsYzMsWJWcrlOPcp0uki+rHnHW9LJkX2zeiQBPwUswV+
/vLqpkuNdHNmLbyD74B5YDA2Qt3TlK2Z82toCNDf8pGzwC/poJlIJo7OPEB0quNGiPs8u+NicDO9
P6zA3dCKjneM+nPgzBf0bDOWcZ/L5Jbje3PDTEhig9AfWvFF8GhkHVxVDD9nDEkUajcN3RnKiZHy
hJLVbDy7QTltie0crxJ7gbloKVOIwYuvmVPGZxDErd+0DM9PuSjXuiV88VGVxKEMFewaHeJbsLp/
EsmB4oVIKO0hAG3jNH5i3H1sMLgKfY4SjRZC2orF5CaFFNihrKmd4oaeI2DMiplUFibBalW8cv+0
TX0V95E2NtGE2t25nRqeoBOgE08XkRVhH1Gtn1EQQxWfbcbkEI3bYlUS5DAldj6mqtZJSJTHqEM6
3N/3bGOtCQZyXBVd34f1gyHrkhBIg1b/epNA6JBlIE0to2Dop42uFY4qH+3fj1lCsqpysa05jq02
qZ+RNKCvgVEt/k+OCdKlALKa6dfQfRDp6ZHQCipUAxWJsTJQgfNslm0HNm/lcrvRFiqU0BEQmNvc
U3v1veQ8XSgH4VzkZjCowzzCmlGLDa4jw9mLuE4fC66dwS+AMPcX/wG/k3IcIk5dO9JpAm559OxY
e0np3M7dX+kprwu7X81ai/W8c3WmMKatdxb22WwEAwn8lUhX++UCuG857kE4HsN4w75lxT7KgPVu
odjnB4/yehGecrHiag5xdRRc9Y4pfut7LV0KbIvcp8Q5CXPZsxi/gPtFOKtfuf2APP91QX+YE78R
yd5G07Evpdd8hQg9TAWi4FzQAosJFHbs3Mceo7nFA1Vbf8dpUFIu4JAU1WQExvg1bOvYONL38eaY
ftwaFiIwPe2uVWGT9lDkZWv1ccpiyodxpt3+syay3K896jg4BHz0slYI8k9vPz6v/xBWeE2q/ebJ
U8QrOhs9UIlJT5qjxOzuA44id52JNlTVNMxZuUcQUsHIR978dQWa8O46jyzkhVObiCMvO78yHf0V
Sa3uMRhwUy1z/XL7sv2OgOI7qvcCQ77z1IBQ1NFWbHzdAn+tOgpUidXA7G9pV4MCWPPTbtpxGFBw
elrX7cfrZR1uB8pROF0/ccYzbPMUwUPU4WrSzzHggS6G//HoPDVO/xm/y0qTKZlCM51mbdDCCgcz
dy9BpeM266MF1U7KkYXu/33x2Bw9sy5w4GINVK0COCtUZsuR1GKbsLUzzilsJuaZbQDYiO9ny2+w
N/1TyfDLvWQ5BSk6AJvRVJgjhhRYyzuL+PBxd5kxlUUmHZNTTC8d6f6quBw8ajB5z3fzuD4rdauH
OAwfpZS+y9G8zQPEx7hUefoVqJxY67/O7JA9h0uEaeUmeE+96pf05ypQF5EoCCrMnk6curu3v1kd
Wt9BcmoBpFGDDVdD2eO2rG8xE1W7donS9w/2LDRNqj2OFKkZU56l2ZD4A6TjS/QKpdYzR8yIgvPc
WMwtrrmvBzyk8v/zQnigybHLnUt8F+4Vsh3fWMvdaLCkRuZe2E4lZDVRZdcXCXIrviJCDzk6GNTI
QkqsR1deUjHfPyS5aq96rlLIvPUqqSPStlSFFC6Ixh0sFYFo7M4Qr4lXPJ60CQjbEzTu6sjOFFgO
8M/dgBV9tLfNW1SDANGZ9okmzhJEtbZxIvwmkYfi/2/tNckYiX+MnuX3b1gyiXZas43Nn1YUFcwO
QihD9yLPCOo7FK5LO5iDq8GpywRUHKO8mzkpmn1B+vQkhVQibs2gB1D5/fVDVzdWmSb6Tw0P/zRH
olYs34eIkpljrkzu4yqGHPsBGYSjMxGlYlGoAaWCA/uuX4TU47ZQyS+gnwsYgkW/8llF0Y+1awF0
n8U3lcj16xyuginiX9PCRJY7vBbVZGjD1eiOfa6D3+wKmdoY7ZH5eURd0KLrLZGfmj7iPIKQCaav
TSecUqkziNP1s+FOO4hG/X5uVBdmg7MbrGFUpLNdTx5vksqEPlXZ37WIrCH2TU5d11yemPj09S8B
qqtyoWk+Uwnh+2uuJp4NKezSHW3r6Yay4xMeycoDQJmZ1r5YqCAAIFW1AVSmF+uGzdlWQbLFFJ2X
GfMuUaPLQiNZxCYvOCj+2WIJfip+I7k3bFSrwgGs3X0Kr+4+njsGe+ncpyIoOWdtjZAfxC+Ov3e8
VFSPKf3vnnFVgW+WIabaA57y/LlBUcv6NF16pWkDIfssHZQGtTiRNoCwQz0+BNJdjW7ZZG2ylpRP
vsvKDptYavBKmFnUpK2zIX5rlLMJU1Tr+zcisASx1ODxmdK9ZgwKqja6s3LfRsb4Y3ZOLjmvX5n3
MHALu4Mx740uyeQV47kUPBJHQuk4onrfG21LTXSb3R/xq+CCCrE9yvVNUS9c8V/ehsghsUURiba7
LSsNTYWIR4h9YTwAHdHwNerslfb1jBW4JtpvBtFB2hOUVZvuTmm9LjlqGHYvL6EkTz8CbDXfukHf
Xk4zNeiYKabsIrX/ik+PVg1X17GvUwZ9OrJsQ0g9Ma6n4snblY+mDXpMSM8EKlTYC+d34GhQlXI3
yXqa0Su1IPED2AFthBlFDxhLED/pDGsyYQMaR8+uTAMFXQKgnKWH3pRc1TJ8DIgMM+TdZsVaO/ll
Wcn0Tdr3DTFgBCgxoZrsR7VOCptQ1eMIqZWeZnmB4fv8SGONO403Fus/I0AUmDrAjJ1iqjDujyqn
0LHNOY1WORKiNI8UQ7WcEBPI9pc88z65HN9oOiMo2M5cRCd4PB2dsjByNbV7X9h6kwJhcCEqePrQ
x4PFrhkpvigN1ghNxJ6rrg6m40CaQaSBcus41xafW1ytitwdAymaLkcWy/0H7I6/iDs2a0g7EN5H
WN+sIu7gR6tXK8swTLQOAavJR4B8rSs93+zgQpfiHgDkcVJJQzcBxsOycjqug5Ec2iUnDJXnWq/r
iKS/vQGeEXZZCYNbd6gPtOgQ7tcSdc7CjtCI4OhsbbntRmWB8IG4bOWPe3uGewpMiW/Zfk3bgBLi
XgliW8mlCsfUUPu3ae/ILc3TJi3o+OcdpLz7vXMo+RU88Ots7u1bjrxTumaP6BM9VRrC6W8NDP73
A/E6m6CMuX32/82m395C/7payWuj6nWsco85HRMrg2yFIwD3zzPzQwwEKO1gtyNtW7yeo1NhD4Y5
8bA29ixQDyN73oirLxekmrSsZX3yaQWAQDTmL2f+5LH25sVbPmK6G0Tf/jXpzWwVQQKkt4qlW0VD
m2uyDr5rDJYVgJDEQqyVkVd/fZabrxI3PX90DNa8KNylxQswRaG4hdGT91Cs4TjFt3jlYUkXayDj
lU8XPpzvRfQLh9+/adlJM119+d6FpudFw22e4tDfLeNGsSofoErewywGVvlUPaGnqyDWXwKV1NmE
66F8rNrUIJo7gBfpV609Ml9xUbtZ3tRnT7iZJlKUHjfYODNRDhc4p93UeT5CZX+8hNLMwwkILC6o
ozC/sE6nj6MG58z4yqmx+LnEFabU3XAmc1O5YW/YxkU8OkOtKB3AiyHrZYfsvzfIm1hoN1L77/Vg
qUpwXceJlpZLUHDNR+B04jBfKDCJs9GrEBRXfZhDYomu9d1saejLcnFkAx22+KTaS2qyZH0yDbZx
Abe6EhqBIvDatDGs0DyOui9iR+V6YyjX0dcYsR8H3JEj2BzKyC+ZbIvwsHimTm3V3ShX6pdQ0wK0
eB9h5XuWEOkOl/yP22inrp8hAhEH0EKhVFup1h8mzSGQL2Xn+1T+VbzlER/e3Mhmsb5KkVTz8CCV
bUqk2HSUr65uE1EoTUKfFKGcEH/Hkcme/QF8eQTHKWSs5IFe5cQla7+jdZk1LUkvbVb4wO+6xfv+
zvEwhH4NbGyNgdOsTbe6lVrr+Siq07Jsu5/2aJ4JjTvBvbuzHd5BTvTIGrwaqqQGtbHk9HcttPM2
DJ5h9ex5AmFQfzPn3Sv/3c6cMTOSoupap6d4FvZwMyIw9STfHupIT90kIiJb3kwC6clNWP+5Yyt7
HZykZkw1cYve3FJv1yFmHuZG22dOvi7FTWvDJy/XAsPPTq6eFU0gOE8K64GuMF0Y/yrGULSPqlcO
FM+g/jaYohr6jw2QAd+QYSCPUBFGT8TXXmlqaMw/k9tP/a9hMKO2Dwo4aRiEui9ORQbQWpmUkFBU
TxWZ3IcECNikjLUMk+RvjAYaZf1obogF7njD5kKs5RYGjOoQ8mTpB7y39Yb416LLYHU/jwCfQ1MC
jtZvSX6Kx8Awo6Rs7SYj+503YsSyMmlzJQsk55870AN7sa5YKOw4MS5Q2QJ8oab9S7lLvt68gyTD
FyT1aK/jnR07rxclqKqS5vfWGHi2UadyBU0rWsoDPLgvkqKaCz08rF6Yb7FGRs0DM4dqsRPthdG9
ehIC3f6T3zZ+ip9lswcJ1M75K0nbOAsThPZEWUaZ5RzWA4W2zOvQlJLPEKYDIZyvGHQx5t2XKs2p
M460WacH2X5vtKPoUmQ/uDyBKOOFHdfIZNnsMoJvam5BWu3zeLG8MOCi5fXPdyA+WbCRmfpy5QlM
FpqvM11uYHk4hnja+6K6It4fKXOXlsBrWoW0+hCaYHO2TByJj9eHLrvjKbFIkd9k7WLnYlhCF36i
lNVCUHeD2iRS4TTNLJx+v82j8cHZc/1oZst8F5TlMHPRuahqHVyz507an2XJ+WIxFmxreMnDKzjU
c7bshCjS7xp1Pd1SqcIy2q4IeMDY0fLQimWIxo0b8PXhDPznGBb/R8R9PeJhOwHilkIOfG8RUxT8
gCX52RaFrEqDJq9die4dJjH+5MFn6cftZB+3V2OWx/kqIBL3Zct7RqhDnKvZAgGr4V/q2SRqk1Pk
LD8NW0K21J0gqZi5D1L456IiDPskm460p3fdU9qoKa1Yd29QeIgO5B3177nU6lqy1BqBgx1rATqF
+voQz5ksH9z3aA/bGYmiCuzHRGaEqhv9EzJ5dfyuN3LTsnAe+bZoo3MDbmms6k4e+C+44LI0k+Gg
OsIoS+N9m+PdMFbw1rdNoFNKaAjyyRGQdzZufYE32VKZrnL8kYthhU8Jht6yEzAtpAp3TQWMl8+n
WGNrKBy9QMH7Jr8zHrSyDgn7BHAfyBnRwtns3V0idobZQGW/3Zcfm0VBGM62qhLp7id80KUFLsdc
CeSyDRsrBp42w1yQCWNZCxcKevxeMuGdpAPVHnQQssc5cr1x6/hbttBWa1mNTFM/rTKFp1GLhWhq
FPq8Fg1BHrr1jtvs+MOGcG63IzshO6f7znOxA72HpqJnFmnyGNFmw5c9a3DIwXDSIGfuXTU1HYef
5rKc6lCUjsz/MTDlkdD2lOA/rSNo4kyNmSCHMOnAVYZAb+u/K/Rt2RpCGD/F9Xa38C0xOWpRTaEs
GXSJ3kD3h0dyoRFfiFaKFbxYK2nWsKyjv6cP6YPOABO/oWNO6HpgJcRroTbFQPgs5GDjel8JLVTT
/ILBzqG25YZBmGehf9gHNEGEDNG0XIPYWG+X0HqozGyOuApnF1ZasL4UGtmuXYEIM/NdUVEGfRv5
/y/KII3BIX8h1Cba58wmNEC+NApXrMt432MDxeh9xpcj8/ytfTr4muAJk65pV2y/FMuaZm8tAt7K
KLK/gfA2oImN6GsOWZIjPW7yIGxLV7fvYwePOTJLRkYQpXZ2Iwr4V8rHZmtWm5HPXQjZYJypOJhB
v6sqi8zWBCdf7v8U3QnTjqGaLP+Hu2f7qbrerb9BBevJa/EkrmoyeVrt/HOLZZO3OJPHvrGsZA4e
8ewIy1+9xUhKDoPgvQ/D2r5hJfxQx+4dOEnrvLyTZ7iv61FTmFd5L7xn7IQ4rH8i3hZpb7p3lv6r
Ht6raGSfze4fR/RvSJ2UsIMt3TkR42rNjROxm1Y7MZRNZ6sj7wE1wEf37VBawn615vMQ/4NlF/cW
JVIK65VtvNk2AIJFljjJ7ikkWe3rpEDDDecObYeKKySs9p3SnON8IaI9e5X3Wohq6WUbPEppIFEq
0+Xjiiyl/ETFDWxU929iigTMYwyM6ikQzkg+cC0vo9P8fmQVfdqhzdUiaM+JKvFhx3DHJJDr/Hmm
1K/1gyClSz9FiHozdf+rhyQaAYSuqoIHc+pKInCNl7hnrnaO/BIfInNkVJ7hBg9OWPAZ/TInl5Hb
emKj/1m/UTyriVT0o1+7HbT4elypubvxUEgblCZVe+6yVV3EpHyMCV+8GokRT3HzgJwP4rgoNzZX
U3bp3DHaSAr/C6ZTjvAdaAnW2tD/s40a0VR/VYEZjfJ4plvQI1sSMMtFihJpo2OaTo8b+JsZXrtd
NgyfZM1Vb2Uc/NHV6stCSwXAspk87wRveSpSKZ1fAJQBer//q5nvTRWtRD9SkhC1wegUL9DE4HN5
GKyVgr8I26g8YDjNAaOgBlyN9gzDhBdARhTW7K00ZVmVJQ5DzqU6m0YVDY+3oF2jF08LDEzxe1S2
0gqCNlhkRMZ+D9p6P0gXfx/WUruxOB1Z0lacJqye7ezD95T3B4ooHRDdDQ7ZNyLpWuoyPiqwL+5H
otI7tFJpp39ke9QykfvwWweMHc1xdrC1hGnAvLHSiQFJ13Hyw7r3mOJk3P/qA5kuLx7BtAAw7XG1
QFD8WTAoEojzWSSeeqEF/neKu5oJjDJv47S/6Oi2T2hzYlA93LjibGm9Q7OJyt9xMYRyp2FLIoJ3
7X8judRb3e2YZ+BYtAi+N282Qh6uJybOAxXqsUEVIRRGeN08DjgqxU0AOi0xWnBFZlFihBpsW6bi
44Gmmj7Oatw/HbsJqWJYDNrjSTsZacmSQvlpXYkrROiHdMJ0Q5zwKHGdmJo9Yybny/HcK+nhcYqT
gCfsIPlBEoDAv3ufXRuU88hf0twGZ10vByInzCaU3TdyFPdBayFm3/d4nfvP0vClF0sAiAac6Z/E
uiGg41zQ9YbhUD0qxJHcUFpAdirxmLzXfuBgpa8h0hQ5dxv6A23wMbLUoAIpXpTsDJeNZnKxAag8
1+aTq7nKUwtpg4YyXmS0jrH7gbRN3urbkTUvxy/124Gm+u52ZyYFIOXwkWgidBFgtRK00vb6LPGG
MDoTE6dMxYqxodvDU+KTy1exy04Fl+GTWk75kI0L7kih8fzis9mjOJfIVUHHed23YaCYIBeR0m59
VtcESsi4twj5PX0hUeJQQQlm+RgGJdQ765vsPsPyfuwM/C5v/w5sgtFEJrcSQDK9/bfPIh4Swbcs
CPNqSAs3qFdAiMcbfJHMgmtCo35a2TaoIL7BYJhDNpnCF/JDsSc24dpwggWw28a6mODPpqgxW5W9
DRGGBuqin/D/F3fW/vIeBIUboMcLu8ilNqLrHGrT75zZGVMO+zikXhvFSbpQUu3HvD/r6nJtTeNP
kJ79PXMeafQ+4p6OYcIZa1vXpp+k7Uh+QK/tiOqyQeqHSb+/YF/kQ2Eq4RUiJjHLMa6zI+ybUmIK
M9MQYz9hInC/A2c2IVgyeO6NBwupdl2nKL/MOjjEt2q5M45de+BmnQyBWbw/7Pfrr0AF2YlaFq25
wW5VTuexnoCERFonaFUGkQzfUybbwG7SxhuOZWDkW4fPvVbqhPnaNgozJOIfYd0SLJnyvxhfge/T
nDq8ZLnN80JaVLe/IWG8vFM7vc0xauipU8OtnVm7d9f9wJMXLslLCKyBpjbDxSyfv2G7BIw190Ib
Zf2sGc6PFtl0X9CfH6vrmgMaBnVCow/wXiQiKjG3gFFZ9zmafzN64KQBjp6TzgEq9iKYS/0N0Cui
vfmvh/6Wqs5JMw95KvJZEGd77HRD1GYjaxYPP+osI6sHi4TUzuIYwB28TyvXk8XMdRgsBB/QueM7
CKOs6RughevY2fCC5HUqsrQW+54p+4M1ZUJMl6p0NxIlPjvOfy/3YXaWbLQXN11KZCyVIdVIsmpX
PBkeUQqKUCcMKh8NJLlZAqoXQ5PXt//eGgRY9oLPYHabp1z1LH/1GHiRy29/T8J44TCxUpWraqgx
OJ/jhC5KasnwwncWMhDgTJPo/V+B7eidbm4AirBchNwXObNArbR3YMkZL1fYx2Q36xSczpZdnx0E
rPxBI8WUhGW2tnN0BipJolHE8hbcLlfYC8CFjxWdePJfzfD7aUZKtlnHLL2wKscNa4eWu5FQ/uBM
n6e7bhhDMNNBMyl5Tfd0eneBNKoqEbPodnaxMrDwROkzpOLhMkDAprREXfh+uXY+OreOgpOGCoKu
VWGM/DqfGJNJfOq553yBlz6sS2rMaQXSoVuMiBZlT3jvisFzNWm5jqg2g0zmSVyT9ZOSfd7Hc0vF
vrOZ3wfcNJUlRjR/uP4qxjB0VanfN7CRDKmBV45o6F8cWdC0ZX/SSQzkMpcY22bR/yqYgWDDd0AQ
M8sWRgYGCCu7oZUAhhFxmKQyWM8oOxOaENVA4gyjJ2j35WhTcMV3PlU1PTVcl5pDf7J5Ti/EqaFm
K/T7/VCmK9AxiMh8EbOEj2VqZbteGfHZJlOwtrp+F1Zaa5P4ywGO7LJpTdxc1qZN/cYZC4ewCrta
Bc1G8LcGbo5qgyELIu3fY4sY3CdCijEwJLoMTng33s5FNyPBnXpUAM7xtlaVXu4xSIY3C7BwdOQE
W0JG+FAZdbEgJ56FCLu2/HFAvK7Y2c4eNSKY/b0gGG6fYupJp66Mu+X3Ev8FgbtQld0lvHgKlp47
30o0xNOT7Owhohm+GIMXkDuiHNbauQH9PsGMTO97JM+0fPB7MwZ2njqBPC4QHuEDaRru2qnpr+wF
Ta5XkwIA+X3ZM85kRiDA5LEr8vUUm6J6254hubwFNUo2ZcX5fNPSpXhN2gEaYjyHSQ9PAUDnTmBY
m6omsGDHmY2iaWhjQWrO9pzfh3P6h+u5zTtfVSWr4xl9guU3rjOgZ6Ac9JnsX9OIMKM05bwuVG6p
9CbmfYa3gbylPdUIk0TLtlbegugNx2SM7Azx4XfziqjMHGqZdTJYZXQfkX1p3OoF1bIAYl1b3wEu
pRlba0/+ufuTFG/CMZtaNaBJPHocf6ESZv2wtIdQxirzDYVW3BZ6xc4GuJgLr8MbbWRXYy68CvkA
ABaOs+WkGu7uGQnCqRD4YB0F41pTe7fRgQEPB4e3uQX2AFwm0PPsX6TD8gJCPYjg6gIaapMbcHc3
c5neuFoYpnadq0UQwvK++iMvhVIYTX0/PEK1u0swA+y2ZHGSFy89pHugim3TCMPJVJKUx7SPN+Nd
tiFXhWlyQNpi+D7eBrwNFm+hp0xPcFiyyuantu5IhQke8ezzubY2AZSmD6ZZeJjYYHGSnFUgInRC
AkZd5zAQQavD+Js9jGTq/aSM2lwMeuCc1OnVdDcr6mj1ODE82oFt6884WWOUUhdv3rUK5urCaFgA
7Th3pQV4NelEE6jd7NTRl5YlWEazrV1SPoREovBh3Q5ev5rrwJi9zgNCdWU2tdy2aeZivJBXiZaS
nj0DZ3AJD7LSD0oLcAso4WDESYCK/wS9/AFGSwdqQ0kH0mWZ0C6NtPaB88XMl0C0IE4LFMhnGxNg
xHAi/04uGwObRxZ9Kje+rYtSpgbWew+wCbFXZT3MkzCImjx9y1ObM0kkmk77SBtfHMVm+9z3wyTR
o68xd2lAW4hB9fhrDWT/WL64vec+KA2cQxuxroENGtgE605ywLPQEPo9ER21asM7YVNk8dDR/wzY
MgCKBFS2QTk/kYsK0Thh5Cl23Dp9MzfU+AOXC7sSawm7zx3IWw0pfoAbo9rqc0Zl7kkiVWQdCMrP
VXR+xVTNLgE24ulwrgvYdXW1gsHtwUxH7KfDYhlfhJXNfmR5GURgGQUG017i2JOyMXm9zYkCx7SQ
5r3DexIUPpY78BfGUq2TjJYv8J2T9wc7PHZM6Av0wCHVU1OsK+VDgnFvmkcJwvZVSHwfBX3lG848
BSnjB/HutpdwA0ynUabB+uhF5JOFx86o52BIdhYBOiTYIN4PYkMd9NKSJYuf9VYDEisz0d5ACGxw
3/Xnf4J+9d811soS97iS3QKGbl3/8DJrQyKjqr6dCjBbdkxoh99kZyuh98PrBw0Nj2L9E5WyYFA4
7/x07jtL3G2m0quQgFkNfi5iw7sEkovCW/3Ypd9HsVR9qGqye9CTGdgEOKK9sUuNDlsh17C16PDz
84kpguWoXMJ+j8gbEJ6lpXT3KaPEPjVuowaf+h3NwwGOUvql8n1Kog7hOzc5qEntkpIsATsEQiAQ
7ca0+Ms69y17EMyph/Wc8eLVTR28vKQrskZU8tuYYAjZPer7MNlqH8LTo3xDVAY3+JpFsaXWWfHJ
BrwwarHqIGokYBf6v4Zbh05zUSb1t4Lbr0EDkE/LPwanO+/4HJfN2T7V/6KQVMI7U74ey3UqelAE
dfJ47onc+kbBzrlMuG4ClOt3H5lNO9tEmJZRfDdmbCixGz8kDjMA3uBiHFlQDSVT79U7KpymrRca
aojRIYmMljtMDlrO4jUntz01cVPhfkFqP4KgtTBjFu7lja1Y/PanYIDGfnUzNfJIGMsUixzhSMg0
BvUr7hC5unsWBL+m/R1MmKgq1i1Al4rYLqw608UIXQdr9lMw1YQX2dLFMgU0IsNTmtZqcR8Phyt4
4n+jgrYBgVN1uAYfChB4PGXLC5uV9zDdnoGdMHwJrH9LRvoeoiIpCqCamaZhylobSMJTJO1XGSGm
HfVwIXYOUE3HBVEV5XmLRG/VMIlTA3faaNzpZueVB9h3fYakgpHE+oSbhl2/n5+yDLSPen7r2bAK
LnnFVDL3pg3POdj9AYnGFgOqMzZ8ymW8Ip7u09ppOF09b2qb+urCp7anJl7kLHmVfH7vuY8zB8Ul
zwtUq+QNsgLpralziVfXOE9QKWDM2NxMIzuTKrArIUbUcBDcalg+gwItke5X1i5NQLBV3drfJULa
WiHij5T4zfEM1D733uztLW2nhcr/ZKaZSQqkDt55iwv2W+Sk0+UPl3hhA0QqQ2c1L4J/wZ/GcIpa
hMuA5RR38Uo6FKed38JTjsoIcIzhYz/TxFYfo9sYddANGGjB2suiSmAEl//hNUOsQ4OM11aRqdNK
1SFDBXWV6ANiu2rebI5CYe6Ol9YsfiMqBA2mbi8XET3PJhuNcWIekOg8doZ3X94lRu8tBpMR6Xbe
jHpYXrMTms0Gymh4PZrNTrEK26wBgpaPA3gh54z+gSkp0//SozB72V5IbXU8Qa7dGCCDBb649lOo
i0V7p3arm/6kxW3aKoBpxawB1qA0DoyDQM1GFToMWe9u6ox6EU6xzqEZhR8U28ACOMm7DW8F0IEq
jzWpDF+rwcqO0ByAc/MuYwdZWXbLD+acxmJ9TQRUhebUDzKPpH2bOlpdeQig9iw3iB9oJmKSeHeN
H6KiMelQIZ4Z54bhw2ykY/thTGoO83izGs6WFhfLkk9arXLyL44Eyf8RLxqPhbC8aVo004aJzCvY
riWJdciQA/RF7FY8KYboFsg8coo4S+hjl1AzwaD6FV1NdGPQfFc/WV2yqwnzFRXN9Lhc3rb/TzCv
+oj8RQNxIZ+F6NhMzDA8jfo9iSTpkc+uM8rrrn4JoJCk5hBYJZw5wYOfKObuPn3E7XP13izJdt+l
p2gM4kEjyeAFxLmRhdOyBocXwmbFfw4nrzujasWxejaDEHx9WE46tgdV2geNFiM8Za0h4lN8+JJK
PX+I1/z/ayavE1EwxIJj0HZujpV7YTRbl2OPfydQQpEBIwNWdRiOk+FAk/61M1eL0/emvJVh1Sve
kyYY4AsjDm2Raek7XwtFwk1n3u3Q183cUH0KxCaDMGC3YbDPgZxCwPNJVhVtXg8uVrZo6Q1ssF63
ZlTg3f/UJowtKe+uZMM9SlckBa8ZB0Y7nHjFkTpGsT0nWU5OPFhbXZnp+4JJ71ZiGAeyE+4sUKeD
DONvI7NChJ1wMdJKTtnAjlyIShsMC9MG66NBAXbt1vtJhs/t4XhZjqVy5U5uvXWNLOPXd2qj24nQ
W3SqL7AMd5T0213ig19HtVcrQ/g9jEcaXOfaKSF3OB09Zz2Oti33FgH2kCCQ272c0UGyja6Q4ucG
sYEKRV0YKBRrI9N5FnEFBchcBnvptlLAD5zmzI1kViw8x2kkE8JLpXa9Mq3B52m0uQdEzFuYqX3W
qmsW5Hiq9l8L/LkwDfpuuVjGKgRaFtQEj6fGHW8378hbqe1RTwR7WEK5gD3xdiExCK8iwFhsep9t
PAlJXrhAq8xtPLgxv3DMDuDY0WEyxloHNY3f8wBaBjvj1dP7eFMry38bgbsn9JUBVO5Xlrj/LCYg
tRJTwlHRCdm4zlKZddM0nZS7hg2ehDsV+RZv1AYyvPk3Ieea95m+3Pnq5YW9d9mrqbsfWh88VLEb
mN3TNulyQCcUcdz/WaCjFSBYa0rSoSMtopejMDnVjDh8iPHojz2258vNajZQXzJ/3nV2cDEiy5Nq
adEJB2+W8uyRvQRV9yoqfKV3BC2akzWH0DlqC9S6fizY+Adiiptb0Hr9azOz/YUteQwES2iMryHT
/jdgcHPNWypmyBxLqyOchWFrgRGYAVgW07AwOjMdvMXRMCxVuLIljk7Svx788/ZU5tuSecGo3XYe
GByLDqIajUXMZO7wTCjVTfW3rbecUrR05uQn/+8fYnVtsajryOnWZ5xr5t2G5JkPXpmm3utb794X
I7Pi3R7FnGNgiBP9oyYCcxdKfrtbjkunryW/rN9UTm7NRPjGBNlpvhf1uVdRIhOf6foHRkZveuFs
3tsE/FaE4qxZd1S8raOZyZvqji/FjYgfFxOJ28VDqS/FUlwOh4NOY1RX/Y51RTi+LCsRtUBXFEKz
8JTbhj0lIXmmhgm7+X7H3zU4MF+1Lyao5wlX6FQxZvbkSO2tybMQxXkHhL1X1YrBuZuBGC5YBtgQ
3+mrzkiwAMl9FM1NDquWFMAy7uR3vuIVM4RzNhiGBBLRigC4Y1Kl5O/WdOtUgru97pmdHG8iDStz
r6OCOr9BFw1x8LsTX5SG3LMB26Wa5VwzBxnLCaPumDtYchx61dfmIR7n1mGKQNX4MBht8QCvwcVn
yOSMhpS77Q+4GtiZq2Es1nO9xzsziMT3MjR1kNNm1x4xq4YrwLuqvgMjjPZnaHabqLUSpI24AdHn
VsUmlV2sj80D/Vf/fSfLDZ0/3ncRV+Oi30XPBVQrP3L8W+bxKrdb94lAdFP1sJ2YRhXvoVAjs503
SAMKXFPJe4+IuLN8nTWs/7x9CHf6fyx2upU97av9WA4mDrzvX5Ab1JVwHDBroWwVA3zDKumOhvF1
CzYFiujTzQR6EYAY7Oq/vgk2znoa+CDTOc4zeEECGUlgAMVmtZA+5cYptVZcL2OIJp3voD3njYno
ItH3IhdsiB80Lwyi7vb8qtuJveAFX/rPrqVNu8leAKqALoLP2uRonw4s/8pADVVqGOO2t+UVuwhb
iHdHN/h/X2BNBe/BxYy6sUDZwbcQAUxJE4Xr9fLu4uzyN+v7rt5ycT7nujRfTjZ/ES9dGqrysMlk
YFl31H6y45F+eZaisyBUUcuxZWTScmQkfgyk0pb6B3XU+Xk0CQDFfYm0dgcYwI2uK6MhjpjTKpLE
77qDF8TuiBgqFkcfAmwI6TIVyL5IQPGLWp/UXI/iuUk4uoWy4ca3Tybud4g11PTHcfWUfwKwY5bm
z/L/UwXiSlTqImDq6zHPUThqPjP0Nk5FiOja6fYcNJtGhWIlp43VTvFCT7BZEftT0wtC2VE03Va+
vWLCVAtrXDDN/UQKSh0t7UD48yl2+1Ql6vef3lXWrzpkQwO1DhzmBl/97FbyBi+voMS/6vUMQ4T0
UwQWkvXZvJ2AuYPha5XNvdAKVlNaphkzNyb4NuephLP4vpiUg5VVIkzN8ax+f14aob0/2rC154NI
EMAvWMxd2HQ59Ka7qn0ZlidGoy4ECdFp2BRNr161Toosth9K9HP7CU+mpC0P2gxzFGs0nIrIe23+
NAJNCgrOY0cm1TVrmAddBuyNEt12VuOYtI/8mAEHtw6sm6wXvOCPXKZI7TobLjIKlqUY1xqlmyzS
jHH6QQWzM42PCWZ62JbhqeLdD34TB18g5tbxmVyCBEq/7lLX8WUoMVoQDDjbeerpxX8sKeIzyvMH
+0mZLkNugFZQn516w3rfmpNdAIkq8KUyJp7YCFAsCGeMd2SSJxxQOD8WuBWj8nL7XcMXWxdY6LPR
MKVefGb/j9fkJqyuSS9wADaK/2Ankbxk1LhOmg+iWJHP8Wc0/9W9Q5n5v1IhJfiFaJERajfE4Ari
j/0kMN7Y2tUh9zw5uzl++cYu1sBX4JJSR6XPH1g8BKjXeuOeRjVEAH3R4jn6f0OPyo4t23MgdJgx
F+MjrNi+/F+I5L+7zhgza7zR1sXB6Jet0pQiGP2cyedupDbUw+0ObmUMb7MyK6GmI+v/Fenbzd+1
f4tBSYCGex+dWJjZF71XEW84mzNyfj2mudQ9qci4OPraBLE/9/LpIRo0lT+U/1ZweUBq+Z8xx//a
NocaxqzIJiOfFLSTjCEapowa/eUJkp7BDVQ+8N4bayGaAT/ebnuBssDXEUFxaktPH+Vwbm2uwhNk
sPZA5/1FJSriDtsw6Hk79QVWqiLRJESvw5N2+OxDKkLzWjT3AlsaW/hGNJoc9t4FL+Ziq0AQzWI3
zG5AmQ9VZO1YqJu5xAgiuJrWcRYEkmkvLprQFNUgXN/WJWPQezO44pFCVZZgJiCP9DBagtMJpAQP
8WTs+Qx6D8ufKU0MgkMgtOPjYLj8xvxssrDjnmh70YqZAQzarwkF+fM1YDpxbaMgNFMqUseQ/XJP
RprmBy12gwYaI/KfAmdQN4zA1LHR3l1Is9Sq9l5A00V0AvQLzRzsXmu/cMwjqHRf6Vi+rbVaGf/c
Ios9f1UvEHgsfA2+6SIgDrWVrtsG58RgWlPsY67yKzKpPbZb4cgAPrdIjlg2buMYo1CBZDlvThEf
fLyE/NS2xu18ITFAOQetxPc4Jn3YE2P+PPlavohFnlRMZdYb9LRWRnEFDhpW2j14n06jRCC+YYI+
LePyMfXGNOSgFB3lH+F3HM7oJ/H+a2XOeXp49vjftszgFAs4rTpgGLwjOI+Flr6ExwMpEuoe7wII
WfC4RAIKv5zW3QHBCWytwFdf5pv5p8cSk7/I+2HVd6tqJAPcCIC06gU9/HqI/rvmSjjGhrYRu0+u
BArRk0Imopo8rDB3eNvIbw4eqwXcYAwX/nElvLptciKwNb3xlw4OI3607hDjjgcG33yYyEL0y2fj
K9BDc43ut3k6MuZqBksqadrML7yfr9OHbcOFGUzw5+IJwdFPXcPpfXEdj2T+gV8UAUOyeiPBLupj
I1sqA5iRBDW6sqE+nG/57xFDBiUuHU9H6T7/AqRpH7iHVJF46Df7bkQaniEotW6SV54BryEbE7yQ
UfhfLoes9AWZaRP41UOSV68GcNgzXnB71NsiItVm/kf2NZRubLFZItjYNnvgse2Sb34UQ/0L7CKA
+irO7KtoUKRrdpT04cP6P10RgbOI3dkQ1f8jTAK2tZ52ZDD57q2F/3wJlctHo40co/oAtl9H+PMv
/JVCFA3QdJrfx/l1ElONRCqlEyiBqgYg0DT+fd56IbIhnv0hSKvSe7h4WM5Kdk3rG+CvDNCMeY/m
jOXaJAN+m7L+d0GWWcNC78BZvU9mvMMWHgHbWhTsOA5a8iE8WDOsKASdFE//J+SBu8ilYbQS6bwj
IK9AC+QRviGmDUmkRGUkE1XoXW/S7KV6RZJ0b7Ga7G0KZbskENXFB9TO2dxsXeA+hDsfqoZtBnW1
kMjY/CTEfC/yvkQkjKAqIUL0r81zmAkfcP72PiYeQoQ14IfG8jbaIKECAd/nF6XSKdw+lprHD2HK
9KCZNnseiQrt6jJwrKVOdO3soj+IfGskeHQ7y9oPiqp8Zwwt++0G5k2ENmjK9mxZXJ6K0hbbxb4s
JyX4TwRs2Bll/oMVI2isOI6bAVV4t9RDxXXrElyHdDNOGB/reU4nDPwcBZSYsg5HfMdGMsHzqJBG
2uRLIk1yAKbUT9+mJVaYT1CCvG+vn2YWWZYkc+nwQqY09Fxo0CCuZ4SyjSDTE98K6Ewihoc7u99P
tSaqVTogPAekhPdK+6XBLieGbSyjW4FADenIKAXtPvqUy5DgFjAJmnkvAuBLAHSi8m4lSOyVWn8G
nucYalxFLzicwU6JScOiDLw+bYJiQXhDRFSCADU44eB+OPQ9u7exmilIU5IpMcrowRk5JL4Kxzqi
RMsWr14kv2uZLgqX5DxQGGCkIkrZVxiGdooRL4Pqn2PKzBb79S1C8omHvz/lntzIRyda3JwiHYTP
l4xR8esex2mYMwa+9T3FyZ9kTSx6DJg9wGNyb5dmX6NDrrJUZTVGFHk+t2YMGuQaAI5y7c/Tsev6
9ZVLLilDAQnrTH6thomLoAX0WqAujp1gkERbaYwlDVtwK8EQSJqOMo8GLDwu5yG56BwWyTdxwpV7
Qqe6eiBkKdkMpz9xHYe/G8KXu5SFdmbqyK0pJ+6eDFIuhUXoRcOULsjUjuQOryQfEfbnu5Eaw1hn
MSSiv0jaD/g3H08vMgUtA92SnlXYITohckyDIJ82RgUDzx5nrhp/J8qM+egHtn16sBZ9U6KNqYob
tmfx/lw5BOQoTRAUHarb3R1/greZkrx/W1SpEupiSdAgSwZ6m3v9jUgcXpJ88Ph0OY2v75rnylzU
n15henwGh+cAsPY0D6sNBla0sLI2UAgH0QKkMRMyssXI8wxSGMKjMYpkDslm16YwoTH2R/hr+LOj
uqEu6nKqj+yg494maCjZMItMBw2Sl3WM5hwaY+gjcaO9unAuir3rpnMllMXrdNXBJHjhwbtqkj/c
BEs7566uaGkEkf6wsHZIS0LsaGy8mTTpiLXdG/Vg5WT6cavVMU0LKG8/i3UtDoWZQjhY3/YCTo7+
7F/1x1O+NX3hR519XtP/3Jcp0oWZMuQfgIiBjzcPobSltKJ+r3dMDfHU4pi6V4TIMlSgNhA4pRC2
6sQ0Nz1gs3ohGAKzrwUTFIXal8cZW90fRNMA4Z4Eiq4kMUBlL4o7Cu1gSCdhbSccJQ4eE/MveVM2
+YMxc44CdAb3K2f6hNxMWHAnzSkTVpLJpb5wstRExhY+Y7GUWxSd98XEQzYnr3V8D+WEqBN8tuBe
6T3S6jalB0FUqPeFM5GYmOPVUbNRmNAeGoN1mGOm2dH3hhzhiDOQEjhumqAVev9MKoWwFuvgOGKw
ENxjPbsJGt4rz0cvfjCegWdGQjT+RvkLDFubhYKFzwgggtdrhMcwUhfIiSGQmOlFGJGsBYT/izYN
cS3aAR32TNrFAe5VzVqlN9Qq6LkkyZ3p4RY7vjT+9ckRtPIz5kOTQYrcj/V0kEDJFfGiu9nYZ4v8
d6gL4R69a7/wPNh1mUlsqVU0bGR3I6DuGBFM2WVw2s7s0hNGKCEnxyyr8sMsXusdajKFWA0G171R
/PslLfpaYfVthjfQu7oBC1nNQO2FBncXXMO5A5yALQjhZpm830iT+8ynXRcVdiBN5iJhz3EOnpRc
AZgwUDnTD+dp2W5/108fVVYzB0whCpgd9HG2iBk8ZHcvzug5HdveUM3JSuhQ8fw7oCzoOnWKugaa
NENTpP0m0A7Z9SfksdDAZrzuLNfalE5qjvy7JFjPH3HgrnIM6Stx4Bcy4QyOn+qqzZJ7zqOLe/1P
H7I4ycHJFUg/c9VGrmSktNZKx1xAbT8s1GQCow3z78TXTni5d85YG8orqUWvQHnCF3uDfjShIdF8
K+pFL2tU7g/FnOB2SDCu5+DYaPO7gIUcfYQ5ree0HGps40h9OUBvwIxpcK3cXGCQ70GQyGXepGy2
/YAR9sG9dfaTWWj7caOxwyX1/v6HhMBXr9xQkGztDGmdD9CVvBGGbKNO27IikX6vFZfCQqVI5bmL
G9KuVkkHDuJvY/oEWcxZ+baCuHseUFMl93nakA4YWS+P8PBu3AfUr9r+8SaNI7sSLICnhV4z3xKe
tqpdz5Y8N8NFbrhYxXSEOhAPhXDfFVclaJ3OEiUxD3odiwxVmV7zTRbd+NWkc9FrQmFxclgTJXmq
xgZzewjuOeG0jLWhkcwHEGvOOqt0SsoCfhnQwosQhgJQI6Y1IXsGdkxxwFk4pQ6+R05ZFvXdGaid
YQI8LFKYKpIGz4SlMXNIuV3/g8+Q+DnOhYf/LNMfxmkImTlt9cc9VyXhMMmShW09xxqeXY9sh77Y
OgURgdiMqhz88zD2bht4m+yijIq0PQOH3MPs+p6ieQ5aJSHDTNdpr0QtkusiZJ8OfjX+aLgewFj3
RfPucS73DhA2eU1eBpekOU2C81bZ+6JN3dGcPw9O+CMs1pqt43DR0noq0IJTCYtm1FWWvKrisoLL
9HMuSf9kqxa7Qb9thk7PpQ9398ij4XbGYPwhPqVoVGT8+dnTU/ZHVrCTQnVGrAuU9PGl+JgIXsM0
7Y+cpKZN2PffpKG73PK0f28odE3bHpZN9OZquO4P3ivTMzygtWP96CKZ/0kV3UH4W2znu3PJvamo
UeJVx6fc1eW9W7wwtr+FpgduCjjSWF47MtfxHRsd8cr7uwAYmhWjHwXqhKcv2j5Vj/2snyXr+2GR
awuvnznhHPMmsa72iu8l+uR0zydQer4iud92qUn0megvTT5Ldw1FZ8LHXy411rLFf5cT1qXPgiTG
hpojA3pH3z1zoZhsWLS2FiziXwpJYxPCMV63pCmC40zAQsjlm8okby2Wn5U3+vrqb2p6Dze8Kh6T
4Xigv7TEYjx20Tmz4ZQx4yY/AH23bLvMV06u4xHOD7693k3N3YSJdfb9AhVwmf14ftsMnd5KjW5I
9yGFYMQcv7Wi7Ypa/vcKtak6BLi3NzxQPTmTZv6P94Gir2xL4uUM6sm7t8kGnayalfsordoh2jIO
VEKpJOWqk6KxD/EotJW4CUt2ueX4h4Uhf2g0k6EBjqzPKBM4S0xlt6lvD+0Jo3/To6NpoW4FP/l0
U2UXDzEWqG0VgtMb3MzrIAwU8C6GiY+YilBpLj5yavth/R4AMdr6ZmbGFgEzWMst3/fDbfHV0XuK
hj/tGK0RRHpuPANbgIFmU6JMCA4Ivp1HYya61OBEuyUSg/N8SKUfJk6z5fNvPJ7zXLKDQuVdxLq/
SrWIN1Zhe4oSallor30vCpplxJ3UrlRS/hvye7p9XAIUfYJgW/NyrgwdAroJ9pE+6zYY6Z+naE5L
RJH8NNAzI7uHICJK/gaHXxOQKd+R/WeLK5wVLGiv9AlgnNtpGgYds/yE32pYtyVlYAJtWNr7i2CZ
Q9tX1jQuXJodVPd0QztjHqatT3FlapHbMRGpIx0rj5b2orfRAZCTFksOKXFl4vq0zpxisnG0L5WJ
oRd3iy4ho82sus5pfjpdO9lmLfkzN5UCLDPUQpo2X5jjXjpFaWKoSYbc3H1ZC1Qg3jgv3rg/+EMx
9Td39nkBxgu1kD8nCS7q2ljNVUz3BZlMbJcpLAtxM10Z4MyF2XH75gsbcnwm4e2Z89r1XRTtXYbS
9xuCvAzbt7nHEtI9YwizPm38EBpsjdYeuDn6vvjq8gszsIFfsYnp70Uo2f0+IzVAGQp42fCMiH5D
dCY0GiXVMiU7LuPuAs3fio6OWYgxcnd3Ufw8wnZCjElfccNBcvJgOR7uM7OERQog0zgby7vfkAkO
hYmGVNx6wgfL5CuHYtMLSYkzvd37Len6MZ+rTSarLkAEZ8A/K+pNNqB2+22v7PgmbU6idT3+4zvH
8S3+8QL7zenkhrn8/fn8871bDPgipsHTsdVnkqW9zRVeY8V8coPLGmvVy9P9C8E5fxdvlvuYa395
agtfbJL62PjbbSoTXi/GKfAF+E1VD7qz4Ejz7RKdARxlyuP+UoLRI5/2uhrsSKHur5CA1b/0N3RU
z66dY4l0EYojPhYJNNXOKQqp0Y0RHAsTJDduv5AROYe7g8ELyCG90as7tXBbyX+V5bUUyMzq2kAJ
5e6C8qG0Ega02OiphxuHmN+EjHjAigmjfpThzJldpKu9tpyyseqhAKzA4oUGpaRAuIgmHqd5prnz
qrhM3wt5Eji9m68aWXM/0XrVfj74Y3yf1RcNSAa3JzZ8Sp+E0AeshA/AMilgqrSuB2IcBZn+dPes
rU19/vOkI+Fg5pFkyLeNszv6q38yDlTeEpDToKtKmhVqdSU+nBVUhpRas82tKynAz33S2VqzE6FA
mL4y0rhc3+eV5EDLYxGAxNpUBVQAXZXGqcqfSpWSMeG3/vZfQUSpTP4xtg/atJopMNwPANKEJGjy
vzs3vJJg2j8xHdxhqqwWzI49KQKEOEw7AU1ztZLOGa5HCc/09AAk2OiCWgDGjx8fSvxRPV+p5IJ+
12jQirKuZJTIYF11fN6krfZjCO/xtNDzJT1kZX7UnuUslzQCpob2ZqB73FMX50fzob1pEsrAvCUH
vIlcumoEBI2UkjfQlDiVJlxsWxmnDG1kTZcFuek8IwuiNeKNURciAQsxKYJWcLUyJ5hRPzhqKruI
nUBbt3SMKKX6sBY62TOvtuvnPDNC2gBegzUNQ8n25MgmTmaMTDap+aTdHjPitPVJXfaQ8Vn9NsmK
6EgiAnNCdP0B3gZME04zrDZoPrCfxrxtQ04H1QCjaS4ZmN6bxwjsNVEMSbU8Ak+GUf9RAFkdRcOd
FZWvHOzWKy4BoBkWu2w7OYzNRBj6uIZ9k5r7OMGP8MnLAuvma/9lkBpoCVSmbVaOcle+wK4P8dpk
3Sb86TboNGIvIPhd6oRz3QvGFINtklyaozicnOvc2pA2MorimVpdoXU5ZsuIX67kToDw/huugd5F
uu/BqWPF/Zafs1Ahx1d/U6T+6BN/ON+TY1Gmw6WpNVSMBs4xzHDTHk/MbommRrHfVf9nD3Roux4+
a6Bt7ZIme5gniuEFTa4zT/HYtfgO05Ky/7X2Jn5CTEP+UK6FN8h80xFFml+bhBG2f+c8KzQRysN7
caoDylFHGI1VpE0tFELkGqx0kuKONIKmHvnh8my8ElQtdIOPClco0MBVcPZm2RA92lPmIam7+ByS
DB5pIwo2T+R4j5TkSuFqi8UOJ3cjywR541Jk6iF8KB3gDuvAs2cg/KQq3/ncIUcviVcujvCHAUee
xGcIdHXdb7omdyP6XFs7ajADQNwnLBY0tD/bwxFY0uA1ouChHomxqH0QskoLRWVfHYyMEKpDWsgr
MUMG6yM3kN6oDtbsSecgrE8YaLmAq35rJOD/SzeyoDrSlI+1BVznVRMeREHISxvU0MYeNfBepJcD
Dhlsx0b2eHxtn+Y8f8AmYOikbnTd8lWpKuo22Ux4BdgZ9fXvntTS0a+Lr9x79eQIv+dsx5mTxrMd
tG3poQYUn/nRWtJ5hKYXAEq9RZ9NxJ4s/70DUUnwmUCKtPSFYS5+fClsns9twRmyp89zTWpT2wFz
uwqVf9gqQhotVgviZnsdvE9PhJ9sdwlz9QaK285U35D5LxOicOBX/i+7Uub+0r3+7hzbd8qqGrDq
0wZcX9uDl1QORwVF9Ec/0jFRFjpfkkcWpdonhAoiRrlacepu+kk+7VpoxySXfen+GyHRrtovkZ6O
yFZd79E1V1wRft+RQPWih2U0obgBCNS0u1/UTvb4JH2ndEINXJdoXfkQV3mU9SuOTReVcT5pI4PP
b3RSFe+C1yLg0keUqveI9up/0yWY+YmgpIuqojQaYZqkgselTuEh2O4GfZPzt6NdBk51sL4ZxGF4
+an59ZvU1ADV5JSjUOqv4yyWPzk9anwGhwTfAK2wDFY5+UAp0yc2wfY2iWEI15fEZhsvLSX/sRpW
43vu6FvtO8edWPn5ohEO7ZE5E0kVKoDjdgF8brLHf/M52/TUlScfmAEDbowb1nzDBFozi+Oo1+JJ
apb5+8vR+AGnft32WBMMri4tSQUKL/ZkuWrJqOj3AM48R3c/0Er4ReLllLyaGxcY8cTdPEBQaLCx
PYSAdN/sdZ51oKg/C4eWXMx8YkJL0RWbTlsHFAwiQq7sS+vKYSoAOPVmijfB68l0PmYxPJNndUHR
fId9qxBkT74Sen0RKvvvnotwsT6xNj21CeRaFutEnOI5BMiKXw0613PyXJ02FZ6BxcapVQUIJFpb
/2q0dQPGOhPBVYfioaQlMt+02hRSRjow9214BsKMAU33+EhOSKBjf5j7iz0jrRxDMlx5y/g+C8Zm
U6iaWBVIfLStnfCgoqkfQfymmQxBmn5QAPuM46B1xiEUdXElO9gbLILorJ35G6crG+P3Q1UuzBGS
Fbsxzv9t78GK46lsd7XKZ+EjZ3ZUWuEFRuTlphh1K0PvIU8M8kJ3Rt8O3NWWd0bPR958HWuAlWzi
VSMixjPecpXUzKY2hdPg7RzGrisse4b3ehyp6ZAQOJTZp95WavcG4EVAzbP2V/7IgJ3nqwerWo6j
FLXeKaB4EnYYyzf/Iz7QFuDGyRv3XnHNusnyiYmiCElP1qdnpue1986gyln6XZRWGQIwDv34zc4i
JpfeAY6mVrEUnCpBZctAT4ozkQ11hy6G40hlYaBt6ezYWQRKm8Zj8YcriI8wZ1ENGxLjbM8EWuLr
/3qyVGOTUGV8rAMS+XD5TvrpZS6+RWTdcWOjkKYNHr2ecuva2dB3CfjjRNxHoHgENnjQeaJhFKNG
hHOxzmt+XrDLOgVpJsAkEV0/7rDkI9jyPMRLlO76Cf1uQkjB7mSB1+tKL0Z04nVRPqWYYZ4iFrkM
LrYg9G6gGvlm0u2RZs32WruLbFKZE00nhpLE+OwKsSWshyMgE1NJ2L1rDNzcoOPNiVZtX/DLfV1u
fh8H0iVbQb7/HsBGVxXQQj9vBGP20uZmaUok1ZebfAJdJ0Vs1tQsyzJrUy/qikrKzZkY6oYhUAeV
5fjXZw5BdZUk302MNz7EnOWETgja6m4+hokAZFEDvwXaz21EcBHYM/oZYfxvVpS6s/T+dLzIzvNJ
xKm6C1+/fg5qWpdGDcSS7MQxcoRE9bAuHgh6SP1CapdG1LVqO4vtdRTUnynW+j6wJ8Y5JdR+5/k2
4fi3XsTlpjH0pGb5FkBsT1CJG00hu0tq14fTUek2YkGJO/LiONUiYNmgkiZVhxqg1ZdElDC3w3ef
4rpS1uyb9uJmEK5Zv2o3rRkAQUwxyv4qL45VMwEOFeflmTMr32Bt5IargW2hvDU9Zz5GNrKYPLjZ
LoDTk+9BRIn0LoOw0Wgr2ET2U7uEj0xMY7po6IhPWTzZ+byYhX9NlyLfPGLimtDRNrIDy4XAcSHe
xPakUmtLj5/QJjVeG+t9AiWGsWWt43AJ+/M4d/I/O/XVYnv3mslxImCPa6WYvtwnEIJehUbgFW41
kGsWa2fayydoIS3Njd7dYcTQNCXcPBB5Hr4AL7vdSE3+5hpaBdOlI73EjwF9VvfFDCJRQ44LAhv2
Gf5m96GlsxX55n+NkADx4+cUXx8IoX6qXTrxcHgX6PvRLZn1h2VTeFN7B67zWMES+W3s7BgeIFGC
uqU5pJXntZuyHp6haz51l3Tj9pjuibZ3S2T+2UrOX/OW0agCDssglenclfhAjxqhavOO2JS2YoFY
An2hV/WzCc960uH/Xzw5JE7Wn8TooTEQYJzYMQshg1miMmjZl0sb8xH19TiRgTpoLBSTPQItQ4Ro
lrGUvRXgkNnPWUQ2LXrAUl9RriLEgiI6FnrNebW0zndYHbWjZbItusQyaBkzTSivp5hOhBVOjzXw
xMdJI4qBbmuxVC8M+oVjPZBqsAO4DEWxr9UmCqIO51GgF2KOs+9K1gh2458wN4tuiJjpJ4R8rpIX
Ho8JPcdx2lPTB3+D5q058EGXfKNmxqQrgJUvWcoG0erEudn+f18U2tM3EuWaFpd3mW8TuWXU2/Zb
kmWRzfccCHwLJGeE9FPYhiap43qfXGUzi39bs1opL7hLu5/hrJnWznqq9CRtfCJAiqdciWd8UBOO
U/cpB9m8pivML9QVs1egdhb3gHJHaZmPBmBEsqvhPmWDxhq/9AXH+IegkuG1KaDJvrjO/o3wZ3TV
q3iCIsysKWoiWgQU9SmfIB3xIhAybDza+bQZ5IeaaioaYKwQtgxT48vwSdSHs9LULs5oYE8BwVIG
9Mi8rEPaRPqse3+uxOLzOqzT/USIRPM65N8FVlBdKYmEXsDvJM6FRFDkx3jzURRmwsPSQVh1EAya
Ze8O8/Z+WkNHcudcVK+o8Cp7taIxwETLNdZdn9rNfZp5YPdO1/Ytf11CHjudCDHBs+wtDXZIaizM
r0Vvesu5xan7fpwMZqG9sXF4ypRJm+hSOrnnY2TskOlGKDKHu0e4gMfwpl9BIsKrbWytzYNByNZ2
J7x2wt3twWuE2vWVxqo1ekyD/RNcMXAhy2WrOFI0xH43mXZUKaAFw3mrWz2xQ6jvJVqAuBjFt+5S
Iw+JPqG0a/Qz8UpjFfU1xzqR5XfyRjcHjIEeNKRcslJWvfuZG/LDJVmIg1LROdAJGW9T5jBlv5R4
I58ih3QACJOO/YaspwmH3KOQ3Bu6TYus4nV5NvZa+sXA0YNnJDmL58tKib32c+jXLGR2Py9WOoP2
Sr7jhSjmnc2LDJcx2oiplrz1zFAO3B9T7PZdnpu4aKr+9sPhR6VhzULr0H0TKsr1xQeWmbVTX/ti
1zGOqVQd4RP/TvVFI6u953TQh0OY97SYH18mJal1iMuLvYYKOA91q0B4DTK4inRUmd0SKd++S+qe
U7K5dS7S0O2D9cyrVfj7gRsYKiRvXS3ptvOadzsEUYahq4Ur3C3vRfViqWvKF2lEWl5By6WP7Ek3
JxE7Uw768wEw5d6HSaFsDyuy7qLs0xg1m6/QWnL2KIRv3JGH+zQ/4YRauU/+RlZfAt2lRUO6amnk
LBGPPnZJw6HyQc6nEAP1nKw6g+MKyyFPSSP75ynxa+W9LFCp1QYYiu4nbIgqPAth1mUZ+rW0qX73
WF5dA0QTeh0FBy0keJ6fzeCM0TRFRbuhbGdxlSYZTrqdYG3fwyKc5uxy5PdI/+26a/stmHHD5YFD
bvZFooJvAep7FulXI4OjCfD5+o65uFRPD8MJftxLv1qV2s66jkbyvXDApwrXPfSjs+CnJjilWxB3
d1ZlNIqelzdZNHCTuvyFuHRL3Bg7ikyYBqPUhhshm4Xyjax02L4PAA+H/+cc6uHHQK6YvE+jZGm9
PlGKmLwM5VUbWlYY6kYBjxp0pa+uLOZqORmWuhiXFXKX1YLY6+ZeNWfimKesZyB6/r8qxPAHdXbL
d+GqU32X784FccTvMKvR2eU5r3MgQaPP8l6eDwuMeDcNZ2M3XPfoSV32p2p4KIPUEjI8CQqa7mnP
Inbum9sOCpFxmNVrt38RzPpn5Z4c0sq/1Vh+YB5EUyXFF3lWm4COXXPtfQvsuXzqXRdLJPf6xT+s
tHp5d1XzWbk0ppHVScqvkxEKH5e9pdSrPs9kWL+/Y7lZ9BcnhP59AYGO7gF1GPYBbcdOel42Cq4f
4vI6YDk6GVuHxG4x0ENbZLpWdhMIJZLKj3wj9u8CXZwc/zboG3SS5wSknn3nGR0VfhDTt5KgH3cE
zhU9Qu1On7G/VSBLspunHIy6yezUxDSIQYfBVCqcG7NId7WKUGuMWmX7/Xjx092hkJXj3PdRbTlY
bdIa9wkDHnphPRsA61kuDs1zjbBgQJd+0gDniLwS9HeeKjQUPZ6XcHY+bD9jiBHoB+h52xlwCc18
kgGzrgVDgFzC/xtev+oq0oE5iD8OMUaody+1rQd/EhB1q5dyCociBmSz2oXsTsZaoXi6oJ19BtIv
j49YEVsxHt2pmafdnXDkS0evqKIhX7uY8/7aoQZkjXCiA6SAIlKtFNNQMqA95s4Snk4tsTo6+wfi
WOnWjn10sMN8w/NhlmIRw2PAvVlJmsy/UPnVbqeeKjONdl0TC4ocwq79/1P7/g9HwRZjkaPhyuew
mHRKL8tWVMEoyWnqMQaUhpRC+FBp2CxoQ00hXTKYvjB86zbQd/gS/RfTnY7QUY5fzvkvevJnPg50
rSyvQ5I+4Hef/1PrJySLS8O610TGQ336NceJ/cog63MjdHdbA69EJJR/PhLzHyFhYGULQnCLI/k+
d3SZhKsnyLW3docgin7RZVa6NgrjXDuM+fCz5inur4SiNXy1DjUeTZSuS9HnduK6vrG56gcruQ4E
dAf9Plj8aWV9h8YO+81IBgHoDXc/rK5A5HKub0nRikXDIQDOvTZDOA0LUeSvIuutFe88myz1InQ/
MByaWL/PZkT5mSNnNO15vrXhkn9EruVHPOskemTUIARz43yWjSGCy21/4DTSMT8ooOtq7WPbqZYL
LbkuGP7HNLQgtpGU77VEPMafog1JGlNX42HLO6bKlvPAgX6kfGXIf258CJQVVakaPevWIFrJngfY
it1hghw84XDKIL4zXF/1Ujg8H0ovuUZ4bIZH4b71m72AOaIoLDZqZ7Je3bX8JwdoDU770hMcD1M7
gga+Ijsr9xLjTPx/rAlQzaGbg1+3JznXCHcWeO80Pfo02lOL/m6dxkDHkIJBwqV0dcclJNrrj1yy
aunmDJhpSOMIfN2Yi3xSFvXv38Xyec3+igLxj43QuxO93XStHgxwR7IxZfFGPAOj34P65mU43hwY
XAzKRfVb+HmVjbBDRSNdS4VLgls7jbyafl0LBQ/t5nNXZnkd89dorgRk7P2shs0fl3zY35cjC+vV
BtkKPyr2XNkD53EtNtGV4G6nY8TKy74VnyFpMPU/dS5zaD1irBrGzxF4zaFlx8P/OAGZxpcxE2nw
QaGEiO08BFZMBl2bxWslWsTzDLyZYGBJu9IuZHvjG593YMbzIY2jWVIJIaJFdC6x2rG3tIh5euUY
IyU1mHmbcy5ShXSMeqml7hGQldAEXuGlL07HBk/jqgcLizPnAyvjOwJ687Bh7y2Ah4dc+tO2dJUB
RV13BNdE58oK6NIJpGys41c0G/OTNKy7hrKK1UbEt9p2wE1LzWJUo2p2S1jPRTn+PQn1+hCj0kj9
JTXVgPZ5bTwZoTx57iym6h0C/3yruJS9y1BTVrjG7E8FWL7PzVtyg49+NXVwG6Wo7tzsfrnAEfhn
8BlgD0u/oP8KtlG9drXWRAE05kR/lIOegQE1buV9g0bhZ95967nfcaq59FU/+9ntnZTWzMyve5+v
MgebrjVTYfUFVn1yjsW7Icn3KGQfp4/VAkanDsenS/DwvnSFt9o6zKcLY/+WfM9tbr9egynIHcPm
w7Ilm8G6rgf+nl2cWo4zajP0/A0eyLmWMch/N18XelDoUfRXbB+7LYRtmkR1/68uZlyIkgBrt1fC
P8QwHmKR/DzxiDMTXZwCo8xfDGMIFSpKo8GJWw2/R5yBEPmII/32T2/u6M+nfTZzzdDp0GZYi+Ph
INQlh3zkAsq9h4vRvweUQFw0fLHtMSxBcuvCY8qKT+TRzSr8grx5aa/nXMuIWfjynmBDcFQzihkr
zw/MBViFYt4rjF1a6AlxKMBp8t+Zwk1i8WTut33bXmZyKs3YrzxfqK4s7ArFAKSshXRlc5MjRzet
T8AKJVF/p9UhTH1o0nOe6DVz2DAS+wEW1x+7wr/9svKbiqCpzYQPZPwPIcXBYIzq7iKjbTaPuH6K
WP3EvWFGIVcBAZ/elKkFsZaVcUGgYUhxDA1wq0v2fLyOVgERNSE1H3A+8Wk3exwEE9c0LJNITlR3
Vn8ofaGy4Q+Qyd8SnEN/s6Q5YFwoQPBxJSQh+NDdelOaQ0DVUQ7F6+4xandAtBaJkNDy/ug22INB
Hzy4XqkVRMtyRW8zWeHe0krpEx0272TE1CEIR8PaClC8HOElNNQBjD/TFNt/1wrvQ2AbmMBknVFq
sHbTEhbZysYrguFGovYxtq0qtGxp41yiLkRvQNck2+FIs0B0pQP53JzsvnJe3nqhA02IINrEBAVY
kuqtgMGhM5ci/cILq8xBiNCg2rX5WT8vlT6Lj7iqi8vn9IVqaCZG9RJItmj1zzTQ4k5CeT2GO88i
nZxVhOkYWn5Ug32R/EPVkLnP8UCLRhH7BlGTYQIc/fgSb8G5IJhm82k51iT47rBhzfTTgDIeeZxh
V7oq6G1Bzh0ob14at0VEw2MX/Rj+UCCB55CoLq2oADLVyLe9GwqWABTkgH2ibRpThO75QOVgjzF/
MPBT1gyDeWGLJ5Sqn5bJax4X2dKsWAtFlYfaaF0Tozk8HE6L3QefzyBTIQDGnxuVCvzkb/pymhJx
PiqoBfTf78pPL1DJ7iMSFVjzpIPyVfBtkjsn8pxxcyRtMe9v+xQpry7b44e2ZA8AghOEII4YWo5Q
nzkJjQK8g1++vydgfLMSMjQbGRhMR2s5M/6bR4II8SrVZpbu5GriYPAOr9an3bL+yO5sxByP+SVs
6rs+xPN8ckmCHG4wVNdvSbq4gCWi6HsguaV3X/llNeZfgQ8qQUZeo1kWghylQfnuhYgICxoCjAli
bCRRxxu0M+9Q6P3PDhnBt6VYTOm5vBfrEm1vZ6N02SKPp7mxsyD/XDtB7EydrELhVJqUaX6ELg7C
Fex57rchPloiC+2M6sfg8BcX56XXaPXG/jkPxfRDksJTjbs6yjgaa1or1Q8Hrs2I1iSu2JUNYP2R
7IeelrGN+hmg5/E/d3z7Cc2hvLrlVhhTEi73/NBHxIm6RmYGNUoQDjyBO6rMnGPiLH1XIv2aA3E/
KIHmmRfaGSstvfnEtwoXq+7z91qf+WPy8QXFUN8jBrAcZVcj+8iUtsUr1lC9g3+CUjvvdsaUIvm+
LgLuN4O5Ezm7OJJjienq7WDtxGeFz2N6C/tEtzDgkS+VfSOaI/8tJMjnal6nPQfmsKFEXB0Rb+Xa
4oMn6xSaj4fPP/Jd1oHbs5fOO+z4FFJ4cyvchYZRIWorfegCb18kr0Rhf5hnyvbfIeEkQHxIder3
ULdedY64/ymGyx+BrABuzIurLmZAPKahsIjYFYllQKMH8pfRU4Fd38S+H83gmdVx69CDrKUceKFu
yVQs6gTMGLbHfakUsWMpyasjbPUEkKASEHDpB7gX8muH9AAOsQFd4ZtNEetFipn+ZgQUz1AepKmj
inHxGAjYpd/NP4fNRtc4WDXwBg49Qw/VU9slbWv5bGkGb5B8XNqQJbWKAatxT04yYZDxCKpKaY84
Enw/0mgb7P948AXn7Td/Trwd0xhvbYKkDJSG7Vk2mBKBqXXqC4IsXE1x6HGf2gaa2vxHdmLo8tNC
F4iznEoDMDD2TxO7e7zeTTRnQRSK8zeCnkq1kNbgfYGxo573x4OWNJryIsMGRwwaubCWPR4eW8JL
3RdNH6kdgjq5NvtlXTeSVfCPnNdV/R8eXM71XrqqvT4a+XFoxmsR095/2illN22jh3uy8SkKiFfE
dlRiL4SdAY16ZteUKb9whI3rBTROukPaSbPbtVWgCWvaP9CUo9GRkTq6qcNSYZe0K/iMAOtlWpwo
f5QHzhvJKgXco1b+HdM4RZzB2C/QdqzTmwlOBtDpwSBn8PPy1nTN5m+DkjEZL48somubVDMSrNX7
bUIOATBT1gc2ggCBiK2wcFhl7cldDOey0XSTLjMy4vUX+oBWCdhwhGAqFqjAbi89FhLBQ/IdbCuY
0KvywyyzWymQedK7EGoG5MF/f+s9aIdzuFodkvRI4sA6bGwR0ytIyLbLAkvyuGuY1i3su/XtYpFC
PbqsGFvqPbmLMwsyy+fL/SxcN1OmvhlbMJllPi3mXcHC8fWVh+Thboz5imc5nLMAf3DCqx0n8khZ
IT4MwBoC31enGP4RiwNfE1djZ4WqClAgKH9Z0xGLAMq4Q7AY7f4uAq6HkV5OpVLwr9y58YdwI6oe
vOjE0U6xyYtkCNwA/0txoJeWUDm8k5b9Z+S1o90Bhwdh+3r9V043PvgTNZ94W8kyd+tT6QHxSYJR
bo6SMM2eimiGtwE7tadX7itfWsd2XEyKd2FjGYsaTHLgDHEOZscfqflwwV+CbTHJ4fET2P72y8z8
aeCozzieq0rY574pEv7ym4S3CZq3wqjXUwYIfPLIULXZXm29BRidFuhDGOPTSr68H0md50Tt8oWR
+AYJKS+96lNYLzsho32RYPw/S/f9E6qw4SpZso45fdXLjx3hfR+n90xe85xhcH3K8af31ZMImpvK
VfgSQpFtAwUC74hljXlGD85C87bvsIMXJpqFDQ3+FvrVOo2xt2rZqyOl/QazEcxPGy915Hd2wMVe
wQgQr4kxVJhxA2wB+qjVU6YdnTv3edR2TLNtGseZ5qYdc0jUP6NWu7PE5UZlsaOu0avY+8If9CGW
vvjUKuZaii1d7h9hW60KWF3OnStJZOQ10KL5AnjlAXOug+MwDmblt9f3AT/ihCrQCV7GJdLiBIHG
LarnCnzg7cHXDpVb5Fs8wBacHHdKECSz8fRsUDamC1jZqyUZkGMiebRhmRFWUUEM0r35daStQY7m
i0HEY9Ip1MLUTr2wgZ4SLWHTL2GmUsjtBygeM1EDp8LadKXg9PC5ToVgbEcV7ajblDlpFUXIM33Y
t9RVxHrNcwSLRQSERRmAiwbtku7nRy/DBq0CB7vO/hOrAw6XrOEKW37/TNv0hg4enfWC/XkCbXPM
h4aPvvUSP31tmD900w5Qp761cJ3gUtfxEVYbltMqX21GyuszHijLDPmBFvGwSevd3vRqPehnZ7YD
GQ7xcBZkBMXz/i+JUx7XGXqPcGcu4g0I16IZVjc03QmoHDoWB4Sg5kgeGPaNmE3zFB8kHCo06E8o
VcwHsr+1eEOAkROR9ICunSDHxj3SmQRPuvGezG+qh7po/hqugKGHe0++JVBrDbMhCrZwE/EUufxO
/JdCnMDABOxIFpx5kl5glwPvbbI6VE8jNwgJXhAEhaURxqFSs5VWdhx6EPdPmH0lWcmO9dIQe8OL
TevpEJCT4GEHkMZrXkdBal8K+mdV4GVS9gIALEjyGexVneVJUyT82+9iK+mziE8glITaLhgttnLd
ypEHqJqDkC4a6ya40rQs4tQkMX4xjtExIKViZHVIFkVCxYvC7x/oMkTHpdywtby9GVSw3GetHG72
QlhhyhCDwx0M1e5IPCrBbmG+Hq2Vyuk6tpgjnSb49fJz0kfc4tnoTErxASpKTjkz1uL07JeMUYZ3
elTpxZQ3a0fSFPUant02axHoA3obH3b4P2xjotxLhn0jEL/fZKX6hSZgKrEaPc8dtG38i/ILZJ9F
dtdJM1bHruSkuzjh9l1UfeLtXWkvkVqVZ4+BmbdpjHXHrJoYqxVyx+OGUR9rBMgPPF+yS0K8kvU5
P2Mb22praMZg3qFIjwrA3EPexa/D0/jwfj3rGRDFn72GyQ30oT/wNH1TpWGUMElI3ngbBm1c/3YZ
F2pobtm8y+SzTy7YzWmCdvbkd6AyyK+E+cRiSACFfTBd/j6qpQRMeBvKtTvqzcveMlnS8wKR4GC5
VLKCT3ZtfJswzm1xdtxQN98NqDWVsNes2dDsKfamDNe9/Ot7E4yOobGnYAhVBtP38j8gyU1f3Vqm
pzJFVdqUChq7t1NdbIgMeYXGrTmyNdVoVxGoPZQbQxKfsj+OQsf6GAUz6XFDvL15Y+stXVejojYL
J2q5NdZ6Yn+QGvNtv7nM7g1Kkbk387TwIRxVJonbgN+t2wbDHB6UVfBWmC0IpRxtpxZlAsFp77yY
p6Dgsiby+Xc0wYK/5Yy/yEod2i7aQbJ8hXYf5BK++vL6nM2QpS4bwv+JseV6lgQUXD62/o3nY3G6
N2AxGbgvxKwLoVjhJCKqBTFYHgbnxeRWDKWryOb7MhWpW7VONDkRLCTICQySz24aNnk8fZB/FXvE
q72R3LLj7+3LTmwnnQcA2R5KHVyYGxtau+WQFv8KXQaCZCM1EKg+7LDkHc15wNfbxvgISU9CIfvG
yhw+g+2UfacIG2CaJbzvmHBoswoVkWz2qiVGuBAnNchUCUtQrlE1KrEkqcbMq9f4QaBB8Ma2eNhB
pOMp22AcsNoCNwsUI1qsyqxT60jJ5/20D7yRPL4pj14R9dvW8w1CHSGKGyuMxVZVom93WYuCn9kp
8pthYlMUbF5tWXipX0XEWS2Pf7enBHXBvJHEY/WyRn9JLKpRKkPCmNcXVqwoN2rSgACjSA+QHXgY
9RmIklGN/2JrtuPVwEdQAg6gK3Hnnc7zW1QQsQMbAIp7onJnIVq+fqK5oTWcdY9d5zj66YVxTDgs
yIoQRg9v80LK0uzYnny3UpjW5inEcUV5fLwaaExH3itCewDMVXvDoUQFyFy+afbl3el15UEfpZBK
/3Xz0N9DvEMKWfdMnoaqyjexebnbP0f9QO6TI5iC1nzfFs88Bnjgi2BGrsUCwjW+l4qEPLFtCfrt
nT+USGgmVcM3AVVCjufEJUoQaaOmZLusfFJUklQjZ7HjDjpZky8lUFgVbFYeBtUoOkHEXmtpJDCd
fDLj3v1Y7fWSiWrTrUeKAIqAe7jB3gXl8Os6X7tHaPWESqt+pqAYaHZPM3tYbK5pQinhlDSPd/21
KSDkR0/LmHfpph7tCwiE+WxTzvdHXhvgKXt5WlT+dHQsaXabDmMzZCC4XXZbxMdJt1uZu0QTIDss
+Eqg2EgH+6Opc7g+BAR2AGCMiEMn8CruWR6qkePCONBzvIOPTyhANDyGZYM8FfuCRQvyjDRfFle8
rqt1+FiWPgV8VlkyJc+gXyFE32l4d2JN6Nh2VSa3HtghY1Ed0OYrhKeAR9vYvyYmhlYjBZwmaLRo
T24RGM8TJfuAfPRLzVk6XnKwBB+uAFWZzfi4eTRst2LuT9rLr9FtGhGDREIbGSFt7TICdfmVsXEC
1Wcwm81o2FdAPHIZZ4Cp99+Uxt1SZ/p+YHnFPQ308BZ3RLl2iSnR5wBXFNpkKDBj28R//W+Fb95x
ajRdwe5ntkGXuH1rFlKrssK9eoXCju/nJZ0+5fkcpw5BsZay2JjzKcjKGefoQIs3aC1aFoK6w5zM
WpwNZlyaVcbccmzOotN8kqRQgrYf4En+giKPuDkVDgCiT4jjPTSg9SYclnyze8FGUF1MyR95AiZg
lJZHunC/GxhJY1QLWsZYGFIRPkqv1LmS8OJh5qqXGXJAXbDaI/0/VX7SpmbRX2Tm5wh929bT+0m9
lB3B3gkyje04M34p3a7IGS9fznh1+QN7K87m7W0o++IEux8h9sI+BauKdFzQ2EWgo1oOcgkQwC8/
zspVh352XONqnzkdu12aC5ubddHzKiGKIcby7rN/b6dDpBpTga49DtzlBDGwtxG7Gh5Rp0hhrEKN
OfgwcKK4mBcwOUc1a3beRSFj9e1eo9GuET4G27zBIGcL2hEsKrnPg0+SAZC4g6WZIcffwEOmXFu/
ZAXo0j4T+mj1qTTzr2FPUHr+fAi/SEdjX/qVAo0pH7xs8ai81qxmBfs3IKwcgLlpYC6r29ZsFTCb
fmUZ3DU2lkidW8hZRMzMtlQ2qFr6RJiD7aXFYoWKD4mz/nVIC1cQ4lCAjljt8IcNLu4kMZgJ2brw
o+zNOfNzxvnHubZhsBqVreLviV8Hm2R7XW7Rfxg8cDSZRK9WAqmdN1iSeoH+o6PGw7/gBWKNYy+V
LD6WT1ZicEeMy+J8OUwjnX3T+KYYoMvNvSGYkqEVRPZHWeND0OJVqQ5WTvFvituKXLP8t9kVB4N4
YlmwdFAQGigctGbFFuMWywJ8QZ6umseIx/XLCmdp6ce3J1AXA4ITaIYD9PGa+rwpK4vV9545Qqr+
dYZ0+WefJU9bK9QmqkSzdxhv10PFzo9N8gS7eCXT0af8bRR2TcDa5IovWD/oTaeb+PPbj36Y7oM4
vIPZdQuMKlEP3DdwRNAsrW0rtE+Czokuh3Cf5dxPWOxjZ5p4sAnNvtUzN/EWy56marfTsO5v0QLW
bokFGKmCAf7YQxDWK37ObmzgasH5c4frA4dhFVrZr1AlQQZIPE/dMleX2tH77MlwQIg5VSk0dTB3
uBMmqZ+ZmbLkVw95J1vbhsSUDjOWafsR61O4DCpRQNypntlfQKX2+QFg0IDT8cCIiRJZYjZzcSxI
dUXuub7VLYMj2Px9LMlo9THqklNm4DDwnWgZjS7ejpKLmS27kOYsjU4/Q1NfSHyO9ra/DgtC9qeA
/G/R1MbquPD42TePwz76TGNNFoYOwrxhVoi8H1ZCthkKnNqpuimqrYHQJqllv6thsgEvIcmBGDSe
HiXrmXeHNxN1mVx5C7+80ezY8O5l6PQxGjcf0HVwc0H7jv2bz/PCg5ywM8TgktIlJSq84O1zAxZU
XEsq9h78MQ4ekQwNeb73qR+g0QuBUj6vq0wT08o5dTnViXd0LE90tORNbPX2hFLAQZ1Mk5NUbak2
zwvlg1nJ+8TOQXUeFAyBKdfIXWktEQQmbhhdrC/nKjmqtQDdCTkJM7Swo6JEuo8HWTZxRvNSydH4
58+CpqYroplTuDvnErqZcrA8MV5W5loOxLCHy28cJ0htoyPSFdg8g+xufINQFRby8v0cclRwgfhG
3hVARCW4higHtD/vEd4DdvvZz+HYuWovKppEu72FesVjAsTYCNRdMDHWSzEG431BFZ/Ynp683am8
ogyF40C0mc8VBXDdc7LTrBlbu1ql9WQUxf7JPAUT+JXUqHE5Ps7zBObUoOcceKUexru2tLOqW6qp
kEB2NX9eympVCDd/VvMI7Jc0ynFKKptR9d3/bmKdR72EGFDXPlwArDsrwVVi8rXyJvb2wujaQ1nA
TTLBN6/4ai+V6ZtAQsru7PC3NLqmbdreYxXrdrzOFOa/nlETx9W2OOyt4geJWbvTShSuxbLUlfGj
/PCRxciuWxV4v37zOszHKaUwVeuaWxvLGq7J5iBTWtsxyMpWoIOj7orK7h/+SPFibt7bG8cWQC30
NK3SyAzkaaNtiHL4kNwaQ1OIejhH5rsx7zZxfKDdvk5MLL6WMQY8Sf3RB8oaDEgAEAbdjSc8V3PE
FLxkTF3GJm+oB2rW8LDBe99+l3AVMWdVNmaXvV0aMr+Aw0rWzmPQjcVNdacSKnRcXr4X+PdTXDvv
iQDI+ovSWow9rQBEJ1z/I0p7iGNwQi1SkCff4Y9pA9p7oXt/vwmCLzk0309wNhtZZYxCrUBnl5s+
gKC+OO7JXk6N/xyItBWaTp76smfIC9rsjO1ysIe3wifhUMRX2oUaJLtYPPiJuLdEQR0fIM4QC9Rh
saS3sP9XH/TG5YD1mKycP8QDuTHmj2QVoX8GK6tR20rJOD2SrPSuAbLWJoAuFisVe99BiOGpKnLg
CZkp8eov1QtRTBtXXV99PUh2JqlO78VjIsHrQzPXLDcPebAh8wcUZVHOIAijENgwLTJPFnLNotlI
u4dOVilZB5q7UbC+Egxs+sPXm8Eyd7DJeQe4k/Dcg3YxmYdobrYWwmeJDOmVlOFrqXM47V9YkXsi
E/V2h5mXgTwsTdaXhvs5ANNxQINwRfTj4NyISPehBdTNqspFSOHdfP29rnBlRgwolIHkJ+rnOX3J
EYo2ueR3q1iABqC9BWm2W0ZQP/fRR7ESMOEXXDr4xQFXJw1bo7K+4mSU2MdmBsg53fvl+exIIWUV
M4H0HrB7AWm17w+xPLusJRFn/XPVZTW+G9fy+HilvVnV/FLMF1PDAFAhhWUthJ67duT9aqULgleP
4G6gSC6sJ+rdZs4SatwvNolwoZ3+nZZLYQB5KHOkiKjU4kBE7hawVIixwtg5mSjAGS/9v1Ze4X7p
+6EQDGvEa1ZF3S4za9CGL6xY9Fvo+gL+rRqzmF827hrCsc6nccutPPagERyzycD7w20wy85CQEO+
iFCZdOPwwTfDwgAFoCT+8eehEJ2pDNIexgJXtJor5o/7c2XaoXLdNx5JuxPeTLwVMVYIMWNl5r5j
CwnT+9XKYsMb1W1ZDZ4zfGmM4lOsj/c6RIfbyJzLGmmgBTgQVH4PcOV5byBXTw6wHKXGgBU/HU2I
nSKvHT5ka7RiclUBN9H8O4QV/I+0YTFzAd7JzAH39QiD5NRFkup506B97z+T8H4/v7OYOt04vGER
kXjmJUUzWTTPyMU8s3AmwE1DOkdLj3TC/QdknhP9iTFW3IwokHoY5JremNJ7ABUhK+AUVpqW9VvH
5DRhMFDtAeUE55DZ3k9FHtEkoKD5cMGP/7sO1CAM/ON1z3blVReTKR3X3ITuXDRln4+K9jOq9a5l
kPnk/hVEu+fNn3qtgHVmO5Y4RubvDViHcivEfouNma0fYbUqN97XFoeXAspvpeL93dZodqPXzCqi
XnQ4cJuiIy266zUsRWnNN2ZwC3dBoJxSZHanU0O5Ky+5PYD63odaF7aYoQu0iL3glbMdbibZLaQq
/Nu8Ny3xurmLVMTZJJ64Xn8BNHaM5exhVnXjZ8KMeVATNFbmRxrelcnXQc85DESceYR72XKrvrtD
8hEZJQhvQMSHn1ghLrpGiT9nL1zoaFpR0MOMVPzhWA4cl1kfMcb/RYqjp7IgBH9jzYpI6Og4VC73
GcM0tcJ7vkcX+cq70CFAIVi587m/s5pZAHLQ/e0Ak8hSZlIl0ASd2+T3BawuZETvlPq4nwAVdvpZ
NjCdmUQlbC5ggZ1dhhZnE0NHdo/kV9voAFueLsmlQ5rBc0sxMKr3FyUlnNsYJaNfJ3ZvfV0lOSLQ
btWOGxvIIe8AagEo4E5YjUBBwkmOVT1lhEilV4CgY6XE9UsXQqAc2qd5EO4XEHHT001L/utRyXPg
nXeODV6TMMVe6inLSxcpUWqVWm4kEWJ9B8PD3VLUeX6MYqWcaV5FTCZu/FDiurbq+BvvxYI6Nijm
SI11FNa/hJLGR0JdLWL7ueTWEauniuVLUby+GDq3YYOm0qsp3PIlarGTcX7UuPCtJhvkSTNoGi2u
sYA1gWONgSlxfCbuUL1rYXz1dHq0kU1Ro/kCgukliLGCHxogZbKV5pNGnimC5gkA4ekDcYNXUC8W
RYHRoAvz1VkugW5riuOEx1DW+a4oAEIrrozub/VmLLPm7uCKjUZ6cZLUXid7BF1LuJUcH3ODs076
41AkxrZ9LavptGsnXcS4+XJnXdmAnRczPPVs9fd43oBnJmhMtftOv3l3uPpwTxJn9rBvYRgrDTfP
eOf6BYJhdhGJADH3E4+LcNA61G2u2f8eGD2pIvwWpOEeC4rf8nkPHtIJh9/FI4ArQGKW3vl7WsUc
1l0G+Q4gzsmUi+bQOTEOOK/g6KoCnAI78uLkebib/CKo3aUY+ZNoB5cPJC+MMB5ncAHUdDszgbeZ
7LWBZz4jg10EwkZ1gs751nEJOerqi8QsuauZwidiDhn100E1opjKa/cYTfynxMVfSGn0Z5x9gz7Y
3PANVFqeflGMHk1AmRwHZQBKhXF/Gy7IlCk0Y1ocHLX55gohVP5Z/rjTEJDNUNMhfcTXsCk82aep
p+yUcrEhdqdQVg2VbuSyAH5ubI4eZcP8+edVc8xv9pddIF7Btx9FU4gerftuL31XUr5Uwot6RQeH
wSyBi+Tz0NW+TycPm87zZw1pJ2BM6a9pYll/F5Dk45k1vUKUUjrFsqrn8JMQSBKrMi+AxsxYpuHS
yj+8KpgRZRlQMkDlJ/4Ll3jhM35lPGOC+IB3/TzfE/PO9BgVEg/m5o9K3rpy9+HFGs1bNkMutWbf
xjwQr0ATtalCIHp4GetkHIc9wgwlRfxi0HJRIJv+2dHhh5feD0KTMPi7897NI/rTbVTbt6kUUm9Z
t8XECeMdDXAQPAwiljrVV6rMetUae75mCbsbdoQDlexF8Zvvtm7slS8mv2tIxLl3HvfyFnvrvKc7
4sB3EnuPv7PoqAFPWwpY4QZ0mILOv/JBSRrfNDY63F0sH+kYYGBDX8ioVPTA6A3QiPX2AncST90C
cjFCjQN0xxbpKpZZ7TiU04E1JTLxph9lN4XxXzL9xgjD4W49PqTMKeTBJmVVkTxNhStfQ49rB38t
J/K7o3De8pJFAx56hW2f53R+gHnT7Dm67/DxGW0hLmOe8GhAJANA1AaetuPv7QUdrodzmo+gUqY2
UHpjW6eaSNNg7goWjUZUu4tjGUFDq79MKF5rFgm30qN/fdPiuBQoAqUfNxdjkpfmsv7UWzz6q4Xv
1nknT4FO9AvZLHcMd4DoQ+L6XENrKERaW8sCW2Kz+fiZ6hAcMK80TlT+tmFWMs0O6G+nLFnO0MVN
5J3LiHDLN6iHDmKT5SxcLXtcjFqO7zyccluZYEk17HYBA54p5ke5cZDjorGcOqxhg30jBtnrZiJe
XMJuSgPfGZYTVXflpCR0d53j4Wrv6bhqVfsoNB/WWFbqDiLzrA0dgvjeEXToBY9TqT53ETHnbvZO
r9Zdg+qdP4s0yyNduKQfysyxGGcFTB2mhVD0G9/DL4xuCZ93RHO2ffYKwNBkU6o1mJPay7++0iw6
9vSec9sYJw+3jJJJAeIOCTHZ4BbNxWjfTvhodIZOf62IVaAkxsmGO/t7qWwce+fJXX0XVZCR0RVf
C0bcRW952m+l1P1bN9p0xLup7M2RnNfbioDOPReVO8hlaxrNe2fVC20U2VdbDaI/3TmVUIoKtQwh
NR9UvZkYRdCaCAQbTHp5oAfV825pk8zq1zAjiF/WIBUSH+jFPr4pLoK7KHbYhrAeLSEwuvsU45mp
+jeFEwnRMyaF8y++2eWKDMtr4aiN5JQzf7Kc6KsBkQCRn83fC+L95RX01YQU6slG3ChnaUo7yHQo
yTeLAdgbcg0N9AwFMR/v3MJuzAIhPqNgBaMLjvznhmP8PNnONOO9H7dPesxF0+GaExXsG7iPBD2b
ZJ8R+4y+CgQTd50zp7bt6fL3ueBcqvMaqKxfszVafo3SeYqoQ2bnzdXaTEkP/4/J3BZJrsJKHVY5
lbqEVt+ccLudbdBU31PZhr+dMisgcWFAwU1o6EWl8/ztWrsYv1C6pVV5as1vHbT0oo+HJONikQ3Y
gtoUtgL0TacGqy2IgzBPY4JnSWacV0POM5Trb9c0g7SE5yWHaPh+mC2SjT+qruGrtsVVka/650d2
ilxaPqk/sQO92JRL+v4McuuEoVigDDv/rCLG09T2AmbCwDzP1xVkIDJ77a4QHZiDmwmoH3JYkVSD
nMlWlxtBFvXwKTGY5yrQTxIrhMMTFDlFhK8EIsGw2FvlMs8PNpsoRR2SFezULRs1rgBh/6T2v1/w
Fdig19QzfwPvXpBo6pZwZD9co9UiSxF2w4OnWR7UzEjzr7pUZ69yPXK4A7fSlgm69JdsM0ohnfja
PT/buldavgRaYlGg+q7TjQx+cjsDF5AACoRc9q+NYHrliLgQQXOrr/mj8O0dsieVPSZRvdPcsG+/
ULy+QHjYGuVIxtmImwNvoOA5blnUZ4Inh8JWtbHxI8tUD9TQn1IrpqrpnQ938r/6CsQ6jcP/Y7/Q
0vjsQTQYtrPUSZmuO/06D6O1yRU++/z2iFF3fH8UgUH+roOSrgslYsjG8VCbgXN2TPs/OQ5hf3yw
vvIN3YadQdUIlJMDDJv0rscziV42VEnR3YmKjSeeeRnwkZdgqD1bB6k5Jo8Xg3SPSCyXim1PxgLi
KX7yu6g6I8v4GWWhwZrJN66g5b9Nxz/s34a8L91As8Gwq6XFtLU97wXT3Fx01Y5anpYsg0Hf3uNu
Hl8hZxMVtpCZzShIlhZJkzrV7vALIzYTmOC20RR8PUZ+iwNDqMJZ05p5mnuEcwu+sxvCNXkmUkMV
tny7/vNzN+UosiCWL7XEikG7QvyS0orpokKDjnSWH7M7PEl3y/s5ZKHTw/YHPaFvMDxJ7AcEhOG0
AKkS5RKRq9+OdEKVVgkjk08Ur8WRZI8P9bgSgCwBLGYHSaHU/ek74ufNvMro0xdVRycWhJINn2Zi
DuVSqXHNCibxRBOplJ3dVrLmdpyL+LAF7yRqDp7qoAuSA4A//zBhWpcYsyN8+we0PEoAqTlO1a0g
tDKqhKVFd/1o8fBuT0Rpf/BPj+wmgtWqIS1YZBO3etzXRtugPPtWycL17mZBQKVgJGADcqevsFIq
83f2xkab005FH79Wprk5gUkDCkhagVRq1WU4bIticAO9s8iRvCqTR28UViRaDTkHA4Xe0/BCf8qq
hJyp7hT/kbVkQ6afS48k/+1I4vJsAmR9bWx3xL5xYp0L5QjZNJTOXnDE87BgBLpzIg1iBxukQ+dO
6z7nXiiLxy/43QrvyJ2uzHioorlXt+gdg/MSg0ivnE8VDad3iy9/gE5KPbY3TZWV2CSDZfVb0zGl
sXRKxOBNJ4MTDxTJLvZCd4/GVUbXz7h3SC5UobZj/eyj1Yt6jZrnzKSZwxc2v7qekSJ/ISpj9L8m
1rigp5p3Y8Rc05923c+bRJbW8bW2tM93UqUsf8etDro/SEA4yirzZzLFTXXY5MebiFcO3S60VTth
NPoomvmTEOam9YTKmWQinAb7sDXssGzHoxqxSBKWSV6eBIIKhAPoe4FQdKNMPP67s3lt/DsrzSZW
5lJix+cd8BAF8WWnE/aujahM/35uh/sYwDChHejpVjVN514r0DbQt6bcUb7inC2T+P1ehkaOjuiS
NSg/zCWfLNCzpohcZW9T0LYj2p56e+DrwJsZamuPZ9RAoK+KwQiYQdi/WJm7QNs/bciK7yq8XJ58
PqopjAfEXqMogAJptka5sv40oKfxn5aJNwDr7/0aMECmcM8iSsB2p55SrescyRnSmhuVP5NScgfy
nf3mufCU2rx8cKkxLmJ0sSx6UR1C+ZEr1EIytYntqHc5XmcJej1g8RzAEZD7Y3uK5W/bqqEg2Ymr
6lAKCxrqcxV9eAiwQrR4LE2+OpUc/e7PdT2kn1sHZT8yggvUKwb6XMURMyc6HBLD3cGROLpUErK6
FLJhpu4Y400azzrjdBX2DIj/Q6k+zJDN01qVSCiIjdXW7qv3Rjbti/VFaLTuIpRaz5qu//uLJsxA
l1kcVtT+vpnYu8wRAmzpDGWv+J92KvILib/POZGtg0HwoJdxOEg8HoLCnO1BSNmWwlmf4saue2xF
BhY4CKFlpwEDaA/0ZNQQwbcDg5xdeYW3eT66QJ0gVn1GwLzU0BXDWhADUHc1Mn7+7JrFTM4Y4Kbo
gqfTIiI1xlRUwsLwi13hrtYuDs/rRQdbnIYButmUhg5gecUr7W6FyhjBXiFLmABStrkHs+12bDua
Np9TDvZ3xGq7NVIdqcm9gwRXMj6CUVzNU22HUYXYkdxm6oUWzI7nQzt53/QgariqSr0oZNofTA6H
uKNfWCd+ABdmeQq7tplg9ZjP20Q9KKuc5C/mVL5sN56zT3UEPqg1QNt/Yw/dr7Km7uSBMoPPrVjY
44nEGrWLeCgbNMd2YjmnZ5tGX34KopuAkfEhDusgcZIPCS4sX1I9YPd+PJlThZIHW44+R6hvUAes
l8etfHiD6PAS83LUV1vWoAdBficaeRgMs/pJwThmIWKwzmVpHkwhEvR6COyUCNAPbBy3JRJx4DHK
s03+Yd9v6dc5ouyFC9nWDVR25G9roa79rqWVPML1frtwUuk4kgNIgpBu7F9/KXL5kS7FhFsM3bxr
OZsYEXB+tWofAFNhQczzFsuZ6S5NRaQyvmWTEnke5J0WEtp85EhAfy0ReUAlu8Y7va/SxUXvaHyT
E0dzG3T0kc6vZ4MEk7uPGlIcdWsL7xptatwxyStjdasZ9V2aZ9kJGFrpF1HhsVKdmDFmUI0JE0gK
yKupV86TM4yKr2IgD+L6jtvPZBWd3ulXr/8YKX65o65DgFnzvt0AfNsID313Bsei/+GbRu3gYIr6
ctIlV0WGJZGCipf+BCva8tUUy/F49Jt08i/BUVG/Xcu1Z4UTf2XSZ01x5LE6MWI2KZhpF7muZV9P
WdslW/XuNJ9LtPBdxZsaJK4to/cjvpP9Ac/NBEpTD4H/Pr/MYr3PeI7gqYb0mqXPT5pHpn2Mz9y6
8veXdd0CDmAuCUWglxaKAyTXEIS8pcplodc/Q6+3c0qg1KmRiyJOmxWOJkYKwpEy1lrWCDEJ7+CL
Tgvyl7VKqBu+i3Tzjua2tQU2GEfK2Ew60Dq36QD7ffCq4YSeDLK4+t5Vyuz09JjxHv3h0j5NYA2c
O5Vyclpz6HY5Eg3NVGsJ5U5hrfTes9wVpMpAyBqdDMg85TeOqSpSjscEni6jUHCTEcOlcEJOujyq
9zD9P8Er82YLqTphzjGmzDhK+FbmnwSxaxT47V3Zn4YnegwbFiLrLTODfmv9+EL8k0idtpsxShIm
adWY3Wj3qUebnhT0NypX+hHqNGewfORTb1NQelHtoe4DaqajnDy1YNSiXzU2UVwlVRKlU7ZyWmzR
u6sprvk40bJo6eBs81t3hABs0lzbT9zFftoEZ/pOV/OapeocgUhFqgfrUKwCKRPV72+wR0/8B6cj
pHtT5yRyDce4RAylQZbrHBb/INKxTrRUOXl0PhcdE33ORt8wpp9ENXEyUgHpRpoxZ80kTaabdBGn
UEg3OQZOJ1xv0kva8FiPlehS5Y4bjDnKEwHGMOAB2F3WpyU2bpRa6dWltyojJj/oBT49qpcW9wxn
hlct5GwpfL4W+gAESUhNFMJXTPfe/XnSSCLv/lf5C2FHPC+lVRv83MXNn7zZs+PYOT63S1csZfL2
XaWg/eckaUIZecCVAvxLUkrlU02GkhtHffYcKzwpQaKifMRG3DGwILM9yJ2aPC+bEgnfgCW2AdCg
Vk108SI07CbOsMQicBhbE39jZs6T1yCPTdAf8HWOUOCsR0qVYFtps/jS3YvQI1k73+q/IaUii9MK
IL5PZ/zJd1Sz3LzayPWUkjhKf158L+YMyEkKrvK90nw1zEiQlaoBCk85d8Kplw1VyoxUNJX7hBvL
MxRItIMcJY3TMbHbJ+P4pBEvBk+67VLREcY6IO6zZ0iu60FZLCwfq1rkD6n9I6iDuLnLzj/UdMHT
mLym5h3NSOnGAKIm04e9IWl1HWf2BgaJ8QU6faIQIqGEGYAej7zjiMpUbSvL6wVLSfz/rC8zb3Q+
Q2W2ozjQ5rUw9TuHFkDeE67cj5gLlV2PPTOGRSmMO1892d4fp1VsY9HjsENJ6Pi7QMyBnuoBnbsl
C3hbhk+sO9to9ocU/7QnMtwQDdJq15Oq63LAp2UYSjSxrmrh4wL1+MnfkoO6poheDRAFp/Rmwu4q
XHXWkR5zY51v83W3frb9HZt9p0ODjv7rt+WE/dSEKQewxabdT1xrZ7iNkzdIE4QK9yXnDw83iF46
I5d39Z27lTUD4pj3rlopBoaEYjrD7WEJaKeaBOTxcQdL5QC/J9Agsh2f9Vw3qrWvdYlAixSXlBHS
x8D8hKGwYfV5pfkBHh3Mdu3wlr8BRwr03rRmzC8r1XdZVPTNlRnar2au2MisGdakBLYOikfPHWN2
9bkRr2grJjbinvWDa65UI41EqhkUmNkzAsFeNVrPSBHPs/o0SKKwMgNwY0wdWrCQkkQu1W4eXv46
HR7MBUw83b+Oh6CS9qaC4DIFG0tSA2H5BUWIr6iEBSNBYxrU41pUxGal5hThkohcN7IltyhBKRil
yywZPileLRdH7gzdrgO/npZkT7qjb9l9/zHki1Yhg/768KHu6BqgU8Rq5s4HEQ5FZ2wCZzspYBaX
68xb1S9diQ4rNYbBLxStSLvpUFZbbfaswo0VQZzr1VcRFidxSVYvz/0nvB0W8JZ1hta3DDYdH6nV
KU9wJOP0nIrnKEkgjm9fxGmpikG5I3RtCcvgC3dgt8k04fVRThRJHotLpYwe8d9SJ52ris/SF7jK
LeKpEXtp6bFzuftclc1UTgNlw2Lbx3KxBLF/cP9N9JP2f5XsZTNR7n0ellxBv5KMCfFn0Nlg5ewh
Un+hy5GKQ9OaNCQKlK/mBh1ZQwT9VlfJX6PcEshpQuPnwqA+x0c3Pj0u2IT/mlAUEQNmGT33jEsV
LYpQ2ADvhvQLIS1jhjyJ2PIH2okB1BvqiggxShf1TL9EZcEFhThYd5i+mAIjjx+IfBHuqJVrU/a9
H5eB46nx10eFZnXSPf3asoGlnE9EcKDvEmEqhaIQnKdMpu3muBN74qqfJ8ZgNfNVJEC2ZIGgoHvp
JMmm1jjlvNMcYSFulyG6hhYUKznDIaP1ZfFd5rspLi7+hYPRxDykrE71FxCCdmwLXYwcUm8duAyx
JMNvpC5+bzjXDPxGz9UIvDD9hVqmh559Xm34S9vCjQTQlHjaF7kKznwvGhq0Q8JS61oAmnpwPYCL
tuBnahXL7EGyqsX6szRcD9FYD9IWRLbfH6BLrxtJOKtTUOkKBK8Uc1u6lXMLv9zRZlIBZII+2avI
rmuyIiZoj8qsKTujjBzPeW3JaAke0T4hsEbmKGvMmlwEuSATtmRoQPSQ2F+1DMo5OAtz1CnBvTRz
ioO4I18Jn4/HyAuNs6q41Z/34kUjg+smFALpJJRDBxR+xKlGu3lbJoxS6y8fTRmBwMqMObDIRXKT
uzCQQVgr2x2eQmibBctoFL7YMFiyjDx1gkLnOVS3GMar5T3EKjyCpflw8toKWan3QI0ICDN15kxm
hu6b9ZfT28usLbXeY9+4Pi+mt5CPuVnLeXEGZJ6GnLBDwpEp1HTJqEfX30XP9k3+iutZ5n49DNzA
IfaT9tvokEZ3sXWKTBTLZwACGRFQBRhqXfb4kqKT749gKJmVjf1uM7OSP1mn5uAov0SGgXEdXbZ2
Kf0cOBvaeVJYGXI1jGG/GyOVsJE+pjvufHkzLLym1kEeseCTGkjWemNUUkczSvLu80GJJt1Gfcw3
2YyNkQHGramiYmrspeVjKvbasX1TBhZR+OR2Mj9nZ8pShpUC9stf5NYF/bkY1dgyNI3sNUOhdV94
U9yqo/mxTg1WrJLP0KG6nb8AiLsA1FTubBEBmF+QKLiOGfe0hxVUfvG+kiOCaFzvA6faar0q1gWA
UbhPdaO+aBjWBiE+PFwN1ZfZFAZ9YslTEBsVvkPaIL3GeuCAPOjJXC7kkOfiFwiBpcE/6Qm3BVFE
tck08yDkrGC0Jw/LqBOe91h4WvA43RsNpK3UZQOrCuyWMGzOp3Lc4GK49fMpxPiXmN54dEVQ3WV1
Qu8NiUTz15Co1ZUmaFMrHFcTcLk1RPxGPzz0JGqIsqKiV62NDlPMuXkLtwN2Pz95D5sx9CKMyCem
Iz9PYaZtb0TPxhD7cvpdoiH2wMLqa1YkKhLLQpSfl2JSDei1Bv0/Uh3IaNBYTsq80EOTqz06EgJh
OFGByo5CEDv6mdZ8FPNs9a02XpZ5UoRiWzVWUPmHW95btviQPCyis02wn12KTzmwW783p6QirHUs
7eEXhK9uk7s5cfrr0mD+31h07A1rzAKKwglJTqwYJH94mzxfyefXoFblkSJ1C6Cy86mbNGvGbBAI
L7Zj5x/rwPY2JqT9FmQpbIfZKarLjgJ6CSa9dArAIVzi/+unAAEPLqBTX4X07jdox9PwEFjV6N0N
g05HMmlCat5JLlFT+FJjc3HVPh/wNLmG0gG2uK+umZhkfXKbj3uXLJwiTlXkpNqRZ6Xeg58iNpAw
h61K5A9aAdO/65yWc3fFYJyfaJZThC4eHvML/RL0QVQEgwnyx0fM/eYWoa41rSmNs8GZ3ZjSVxG1
Fhq9v9eKAajte4sN20ikVe8D2mZUrgJgW49trmRYQsrLIAwcO1646t5tDddDzvD1b7RwNHI4v5zW
RVSunv4UPSvD+2us1YykfcYD5HoDcAyXyhO0QjITE4SV0Nwwb2GgWQcklrkoQmiFlQWsIIQAu7EN
WRietK884/WhSyP0Fr5SXZJH/VTSzKwJx3t6afWlBwuZleHgRY8Mk/khMX1sGxYmIaDFHcJfTkVC
6sVTrX6v7R0fto5HdC+JRBjxVZn8rvERTxvLY/KnKhMZ3Q/i2wxf3C3LnLXME3ySUQqujhYGLG62
tUduRpmhml5xCcM+qfV35L/uRZzu6g/17ScJijJer/MJFtKqUfTmMRcg8ctKdw6bJ3W3GhlgpQ7y
O6iHjdeOwK7XHT50xzwBxh69pIBh2yRN/Z/SEPbHoBygh7UHMAFFL2Gk1pMlm9Iw4WRoouNGvCXy
ytZSUvG2gNfkuKFsyZxQfPXcq2PuGElDMlkOCwe8Czgb8QwUuYxJ3ad51Qfi3AlRpxbvtG0wWyt4
7YeZQzDZ2JJvMKUzPTWkTMSBKx0FWV8vkiejHHvu8ps+ligCwUvod6YRdHFBe3pAZ6RoQ1SVZWFS
F9zGCb4JHBuj4VWUjPvtJjgivZ+BThwfO0Xx/iRhfs8NVOlr7LA6uQnhjmaX6ROhmfaDrE+G9soh
wZOG1WNboRj4JDP0WidFam/bcyD/LA7Md+fDtS8Ar8IqksNJ3A6or4SGlYGPD2Z7itvm/q0QrXw1
zdI+f/qNrkndrYDarQvIYocICTGRLd3laMpuvlNiahvxsdufx9Ked+cjcX1RlaNbCR7KNhNY//rz
czubUjJQqcjOWUuz81J5Dw/EIMfjHkuKcdUOCWthD4ppR05nO4mNIniusEU1S8Mb4WpieC/WG37j
DMhCGCOEaAXrAajewI4w/eBWKFamnGbgdqb0ziSe/GSQCj9sDYCXffpPLF0B2SAIDR12HJONIGUp
ukwl1YxzFwKEPMhtT04+mUxUjUf+Gz2C58BkS12OIdJyENnjHo60wUpGVn7BMg6rMVDo3iVYZ6C1
mHWKRkkLjqR0wTTnHad5pRBciWzUzAUuqyKeMWPLxkYIMGkC/BHR4QCtNDUAd5hx+wlQZD+Tu2XC
SEBrn7CXUi8dT9fFplEPjUxsLSaEJhJGmEdc0StTbKozHwoQDCGYzEn8zLLhEdYdISTNnft14k5W
up5vO5yNucibY6bJZRrLxPqF9b1GCadeJODmSdFlfJoDwZELnp5oI3BC50Qwz2qTEo0upwAZkG4t
lZ5raxvMgllE6p8cfMi1NSI72N7ZwN90QdQydJcti9p6f8lPdeqcDIgfKSfgn/0Op6PEHMCRE2n3
KN5v8hoEYnEHSunC6hH7rlIF281RKY3OL0lrralU681v9OSuG1wVrkDWIpGS96/ZWQ0IKV3Z04/I
d1Ofd8RYgqa3ULgEaQE8jcJnEYtXxh9Ys6oCLxdMuJTcoiGaCf72eYG/TbeOYaEc/nDe6qd8IVo/
3fvsCO+vxfcH3AazRWG4YpHhzpGZzKs+Cu6zOkS0eZRpQj1k2zuzarXVDCYDPFM2F3gFZA9GaokQ
Gim3jc0GjD8pcBoKNb6uWDOyiI1GhJhF5ikcAfK/c3ZFWu1jwHoxwduoim9uCZolwOROhXn5r+jI
tLZfPKWM5PBgrGWTD/QjN7pRd5A5/48busJnDgOkkHL0fn2r2zWw1YQ6MOsRA9cSIoNNxI3y9DJk
7g0z4C4ElS1MU0C0ya16bIlVPNvgoYXHvBv9eSSIUYjr3Mz2cwTY8nv8Kd3luiZ9oxJNNpOi36Dq
18iYW2Sr/93naWPnIhinDTfHMC84Za2D4H6YjVoxXWn0kupZr7FSNz2pJ0MNYC5+ncsXI1Zb6aLU
nqZNVQP5fdGNjeVIARFx7b/JOAim0LGpNEc7hE32byV+l/VD5stjgN7S5KrbKnpfqW4iCYTiSatJ
/1B37DoFVKP1Bo02VeGHw1MUakJKpguKlt4qhdfstTWsTZSyvLoAnIPzQJlkvTu8wmP4BlCByaeL
ogACPAvMFYDfM1rjPAv5Q0NTcsQY7XbNJ/XZsyIK8Gtavdu+oE7JIQs1Rl5zgr4aZUpitBq/666V
JTpIdGfFOwvOwoeVl/uvzg4y5lVFCbPy4/okBQ7eW1HKNWxc1MwK9hbtKjDqDMHOcQU2bqyk/KeI
qNHu4eJB/iFi8dilAmI84Zxq1Zs/kaeouPnwwpNVhXYIpyCbE0XOkBXhSYYisLtiWRdF2RpQuJif
kZhzZ9Rz+abHzzQi1Mat+v8ERKF+9v3k2+Rp92VEUP3eFp402UbQO9IjQlJdQqW3Dufkg4Ux4pR1
NFzotEKHpTdy2i3WE5uyfg+F54YxNIo9PFzFRdXZFJvRsOsPT2DwyJzzksXQQpy9dqNuUxa60uTa
dGnvSjs6XAMV+6eav2F06eKY2zx3IHLlE1TF4Bp/fQ9b6uJFyzqN+zAGGI8JsNIEt9z4TI3w/y/N
kEnBCAI1ugbT4I8i3zHDCsayBbYI8XeTPQacq6jrI8AUxlLrEJuRt/wo0MDOuJZGfe4XoWbw/Vib
uOvdQaGcaeq7L1iw90m4TykWpi8+0oE4j5StILRMhPmqoufQxfGvjvjX9/nOdCSLgb0rVyXadfZK
K0xY7rAFSFyxt91vJl1vRll+Z0H/5q5GF6jvLyX7bat6cgccPz8Gr8HM3ABjAFyio18OoYw3QBTd
K/day1b0v/ZUBdOyP+mHH1fF5pdcH3HFg01mFn61t8JxYxZ0aaDgLZ2uMJh29bmqA9tvuR5Fngj3
gRN0rE1qHNi28FoZkUQkDvM5KzUiQBrJGI5f4VjEygG+DhRK8Y7ICkgNnusnTyysE+ROk+QLoyIA
3huH0J9o8L2yRI+ylEYW2foYTZD7YB+KX+u38IhcnndNfHilubajr3nTuNkIIFCpk8AwhCboJkt/
00mctjaGF5d05ktO+1GJqdwos65yBFCeZzjkVexl8mh1h8wVFB4uKzv0r5uL8Y2c0J07uIo3cDOY
poFitHyytqds+94xzMV25gM5BaFtw6KqzOxpR1Lg0XotZ2U9WP32Kd7p0j8+BYVD8lMa5h+IwZbp
a3BzJa4sKiiA5R7ftVdl9jmGTD6/8r148Zgl2FLODjV9qY5yTiPO6htJoCXRDwsmTF6i7doKleP4
tNLWMC1WfhJ8maI+KVMKogwjWoafkkWUkgkar04rvatlhujejzy3tryXnom0UtAwTJR4q+y8aGDT
IywOUCkhCEVZkUnK5CU/3C0ZO6XBzs619PI782mzGOyDNrebcJJpfXWufb/Cl9DdxRTQEdOzC81J
s51ktihII2JpI1FsQ07N/h6rGdGgX1TmT1LuI/wMQblsyOts/R4jTBz9x08pbLVOGbZGroM5CNIa
XgWMMM1yhiWB4YHZA7PAKvSVyzozueysmVnQpwaD99WYYWR7i8IeGeKw4/n402BfCAiKWk+S0paL
ps6p8bqSZfHT9QdoyopYGuI6m1OQoeOAUXhFn+fPZOqvG2GdHBAognYsfNg9zVlgoRtFWVZ5kn5b
+IaBQyYmPFvTMRZMeEaf7q5wQcJ4YqpxTQ6vPv8KlAmciBR84LqiJbGPG1YQp0sQi4J35U22T+gu
e0aA/HHeSMgagtOwH7hUsQ8/scagZbyOGkWlc7DCIinq7iuUOTNXohIoVC79GhEBaC9A2WdeDpSr
ZNDCZCEYFMrWrz595ud0kwp0hPnId2f+L3Ckhyj3yoVm1NJY7H4VZboVMCCcWygM5M+VvTyadyLI
AJeJ4TDLakBJ2yQNjSHG5n4vcq+6ELqSX9/uirG3sWdeZTAsBQoG9i3IKvkTJA4gkhIS+kFpUl69
vpIbf1yga+qV+SbABRYYsEvGl8zWwFV70/xdYGdSJdgNuUNNmnJnnLsSFVQx9RRv3u5E1ijxBFNR
w65yWN62yTQZ3svOVcp0A+eP2dSBRPzU3XKoUzI3uNIKLBivg1Ibhdr0CxJRFErQPFsJIXU2vwGp
BqPt0GiBuj8Y3IN+h8+nSt1ARNiKyia23XUUxWAoLNbUoHs7zVOb9oP2YaNaA6HleVhoxPrIboqP
6uI2uOy19AyVxEJcZDYHbOFOw2KHvSHqQ1rwWy4kbjVfCIoy8J40Q3iviXZf/v+oroIa5IR/9bri
1LWhB/WudALIGsE+PXTPHNf/Fk9Kp2D4nhVeyDa5I1guXkOfH1M4XZOApLkZKOvEcx5KpRAigdoL
8vg5y3H168EwXL+uQtyHHBLJo0wCkm7rAgGON9QvY8jVANWsOs+EcceBlF25+HwNiRzpM+opt1gO
qPkuP6jWH66cgs1WyAVHI99sP4mElaQ3NiWPGkBhQMpcFEzdiyFnamX4Qi0Qxtj+NumiLuZopXL4
1AtraPXQlDvgU8mBkBvf5BMY4tf6uba/nW4HkQp28PbYREHSZeXam/QjL/GHd+0jpRhDmwQeFEEn
RUlkgmOo+AF+FOE5lU6F9KnCvRAab+NmVUjN2hm+BrWOXRxkA/f6M32+H5TO5o3BWgyOebqrCVDU
SM2uE+I6nkcdF5pMhWN4jvIIG4QeBPmc+pilE5tmZ1nLQXML8plui4lnbbtMm1KCHYwFJtWTiKLX
GBnF8g3Utv96XnHKbaR+LDjpjTeS89bJS06LFIFQLlIk6cVp2Z3BQCaziCIKqz10cPxlXP08ufFD
gZDBMvko2OtIB+GETzGFAnVvSxHR66Dc9Sjiu1W79CmKG0FtKx7SHO6d8dBVSsXwWN809/ilLk9l
wmQPDxJyYrTEkkwiBw6e3Mp9N0Tq/JGVYCc2IIGv0fE9wK+ZE1fXmplJiGr2fkLIvdc6R9TqslUM
YJjsFWnspXxLlKvVuh3dKj4rhGno4T7XDmUlgPPAChhu2WKhdHYoa4/1dsm8Kmn4su/Bpqlg5VIA
3/JDZex3Rlx/NtVJ/W/xJVDI5ynmW5wYM6VBZfNgL1O/OQG7dBu4125Cymgr3J7M/cchvtuO3cgI
SF90DjLchmlEJM3fUIBr/mNAac+m79ohHdtTf9KqcJwSeNqf84T7NW6zp3I08+wvqYUM/eGn4Wip
qsroffiX65ABLi9G+ArIz/6XtRmlEwE/lJROHGdWSsUvadiLPi4YFcUYsvv77ZcxExHIG/NAlUZy
Kw0g/Cvy+/Xk7MHEU2cLliG9hGNe7k42G0c8TpHrxuXCQ7tL9Ahge0/p1IK0FtaelFbuW3JyU/7K
G+pQPGMpGfqz0OEKwW1rFkk2O11yNvwiRuasP63F4mRKQZFzbZS5IRWgVtTUv+GP1Mrws2t+B/iC
mhmtp6e5GrxsCCItJA1PSHVXF5FVU5jpXIJoi1H5aDdZSGQKfIyU+xdnLUFdvF8JqKIDMpwYD2H0
xgJLVWe7tU1KddsFHda3hnmzuzw+7St8bKhPDzH+pwQv7QwGg902MkLegjgwa4ICUFwBVRjIP8It
PhdoRyNV6NkNK8KjB+7vGVSgdlZlNcp/g6bmwG3z7uqHLmPljuF52aaJsMbYyITUIN/9UYYTXqT6
8Dg7q6ZuoVBG1CX/y6XX8fbfH13YKJC7SDTvSzasXvzOK3mSOdbF2x02EjM68KCfmnumIZW86Dar
CBrw/nIG8tU1n9k4AFdv8ltsDHrCaomP8YK9X+XM6+Cu2A9FVwzcdTsSWYJcb0P4Wuh/+niV3AMc
KqDuSY+87BMjDK7Wn98J6Z6D2/sL4BzoOGXRjhEeXqLVqbRaktmiMSVPQvgPjxUrYOZkkikfwPWT
WjAEh/xIk3eB5b0bpBTSQum19FlIk+uxpAwxs4x9U8WbPXiiSOYTY+mWwIT9d+mAt3S7dKm3GsYu
ZzTylVVRDLWauqIi+7uSFQwpmlbjYUcsQy1nxHxLEKNZa5rOoKMRLhpQCPHrbtDyYOnr5CGf6Ve/
mWHg+NXd7onJ2mtBIthnTWyoc0HyzNe6Y5UwCHRlE/qHO8M/7fiRJpe72XTPi/Lagsm8PdcO776Q
rRGxRRfRCGUIbjA7FgRGRtk0tPmLt4H/mN5lUReU9bkmhYRsVTG46fmZjXWOfIr1rzaX6jBXIHRC
ZabUaBJOPfQWRvOmn5YmRQggOdgd1F0Um44vFj9QFTSmZg1KkuBzQxIFh2AhTAXLjfMq04yDF/Gs
NYvGVL5u9yYH9HWStMCSL+amAhVx7eoe/VoK6WSz37hgW4Sj027/tXjnRhz5Oh5FM9rCb+jdQIL6
xUQDuZyJ10osu7DXomivJsKuT0pmTytDb9YXx661buZc0+G/7ZiUeNWpEN7Mb3xv5HppxLSvpU2/
G0oD+q40ypipXc3VY8fEw9W1TnduvOlHEbwN+oF1xG1IxgICrVT+WwFNIGOCTD9DG+W/VB4iqWsN
/aLUiMi71NlKA8XRBE8Qb0lGC9AOCd+bcegYUyvgUKnbjm0X1RuSzBsgTpaFf+yooDJO7h4hnqrn
V5O+czbx7Y1qGI8jZm3CfiNLgUerWYihIv1LGV8y+dyMg6owkHr7OoZTcZ6VW/GT4HZDLplxe63k
k8ByhOy36mqBXXOpMRmytzKVblZq2BjlxZ49UD1jho+ND7JZHEe6VeWAmTRgsWnbHNd/APFMJlXv
Z/mXXQlzqz8LVzRYlibR2AtvdWoLbgfManaq0GMjCIjGiUL/BwNkShbNDEED+alGWld+Lu75ooAO
CAEKLaWa3rM7DukcKgMAGLvhmANvf7nktcRVVkGJ0UrYFq0rc+RL8zyStCWEtD62uXdm9M3NM8oZ
NVXhAJeSS8KwiT85Y5kcVyS9ATMN/PohlZz/2RKtvgRwM/RZnTER3a6bynMxmKxprFmI37w04Dn0
Gbkxhy/c8GR86bIX+RNfQHhX2IV00QZQlpzfKyGQGQzcSku2SUvTbLYuYZM4HIszP6lXE5xZJaQ7
oNza2yGzOkprgltU1HSxVO0sd570JtHpfvUMP9nB0VaD8A5BQ8AeLVY9C9rDAVHVGpYFKsOs/8mN
0AVzQzT2C1Rghxqg+3EQ0bpSJ93+8o8H1XqvyMVNwCfErzcetpHxRsNVPhReDWUq0lq4wIWsbCbH
Y4CQ0Wf3719LDZKk8mYS+YudKToBskSLwe68v+VTcT9AYSmyKXiKV19NZSc2DahSPve7jEt+53FF
BFa7cUMrhIjpov1wcDe70XvwGWH0/KaEs0TYi3Ke0MzV6JAAm+CGdRPS3tosR0OO26D1OvXKoKgl
2jhDNszL4Ra/w6Ko7PAauLGVXBg/eBkdAPQfMEkaMnKLQ37ymsmx4wG9/CG7Jh1z0b5E7gG3WP1j
LsaU8ugsEEP/pFQINoLQ3ysrvJfH9UJvQsI/6dwHhBnQB/MKsOx8YMum/VJC8VuNOpdVZo0RKnA3
Q+vFyiYxODgIzSXI/71vmS1JJJ9MAq0FCoiCvVxPkH9F5G9HRy0aNfcWNpvsTTSSFEUw3Dpszf77
xPRAgpSIbP3cCGQ0sxWwX3RJE0yvnNMdQQy7n3ml1nVCKejkN8wdoqtPi6C/AKrM+55ASZobewZS
YCQiv6nIGdXozB79n0XY+3s4wph8LVZmGdp0XE1xTgUju/PDZe/8gPo8jAUWSCv7Hmbu7wJ5Tr1D
/23thqzrHV+8NfU/jEaARM/83Ic/HlmM4mgxIWDWgQBT+IrsBExRUhSQrlyAeIhfFKZ7AxMc+GwQ
HOBgSQ7f1VabgATTHXWzDU6H6JfAoBbSZkz+Uj+vpTWVGQUzHNcv0Ij6mpD5WsocKI+TUTGr3i4k
1DrF1BbAotERGlJ3cd3gA7hlWl7DewuebdgljofwrrN+wji/UbaPq7woGbVnXP6ku7NXDMAq7ZKZ
W2kJNofkw1wRed/UjImi8zeyWpnQlaiMj8dIx9NqGrlSIdqWy0fHnmCQLYam6bwfOZvE4HIlkh80
GFRYZFPHmMo9omvoE42J0T8t3cYBITBPOar0wUbHFvffqKzqA1x4o2Biff8FHKgI2F0uhlBhBCJM
2d4f9dMYhVfYKqR/hajaqZ2QBOOYGH8bw3rilYlQjwPa9La35vrMJ4LRIaAQhroDB50xl3IIHzwy
FGr4cQQrYMntecEBhldsFiSByPMRBYe9H3F6rnOB24cYhGOwJZ4PCHntR9y+qGDd9bsxoaRtAIje
prFoHdNZHQWRmhMiGcxvlXEWzej1JZFtrsOOAgZGc/rzBmCHoIaP1WXqd2tSBs7lpWOEcAVWI1PR
HtjFwueg0nOt4wkn72pJc79+tIf/pGVtKLCWkj5/E+9YMdzvh0uz2N5m71xEiig24uUHbEYM9twf
Km9ZfGxUplJ4L12E+Vl5JL6S2yWJgkAHTzVi3Bo58madZZm9sL4Akkn2fiO/EqI/NI+2e8rilbnT
jquzbXiplnVCcZ/X+a5yr/mAACrCZy2WmNEi0efQwY1Kcj8rZDcPH0urB9fsg3J6xZQPq4gDnVT8
M1oBKUN3ymzNUyCe2EKoVsXV9FyPcSbS+xG7oc/IFgMewoEXGPuCYn3/x10AX5OZHI2aACo9wVEl
wUg5vVwppvZ+i6Ooto+G/PTPEsqPVEZERqk2eEQyTnHTAMLKLn/ht7IxK5bQQMSRFvvQcMFuSE6U
2UdTBOGQa5Az4wk1zSHvnsJUI/txyseBkXwvD6al3HBKGLf8RXLfS+L25Ux8/qyYV5Op3TjU8/Eg
K8G1dBSMtj4loNb+jpPTqYoDE6G58kRsrpZdR/Pa9Cd20gz+vnQq8i+2xwNDuAB8ZI0iaTVf7dJo
Mngt/AzlqpAh8ewG2Mt5RMBz06mwLEi0RnICYP8m2fRjVb1u8TV4BpAGuh+Hz0JpWZlnipvx5r58
mjRxc7Ls7+TppCMcvILEQD8Jh+Ptnv1u8z9Qz95UCKRjipqTvgPjx9KSAqe3xvCuk7df5Ye+xmW0
71g7quRwbRCTBLYbCUlH5p+8F4TSpd6VJjjWG40nK3YC2W5u/81Wg+qQPQpGb+H6DQ47vnlsmkkd
uJuPK2ifHNSLKKNXHlUvcX1Ec/sgw11XTHAeLsa+Qdqpx3NxyXoKZJBuvXFXm10yP8G4l0OLywSm
t2Vq/W53GpynyhVPKr0gqGNgrMnMIhabdNcemgyMFI3FhT9j/bYNv8yny2KkiuhH2MgZs81eI8MI
9/gYGWeAvuUpz6k/gW2glYzLfOEHS6GPiRaMjwDWni1jXaL018OMaUmdQBBg8LGPqo2DkwhFOZws
01VqBJmG75Mos+ygOJS+tQIJ8K3aG1xlH99l8ffYRYyOmerhx3f9Vr/XzM0Nqz7XstJdRq1QEbGM
9hwhNPJj8RtUeWneZTqdn0LaTuSRNGy1hZherh+vlA404L1gJyJDDsU/teDosqfL1Dujsu+C8vsC
AUO1mgLwM7LIo6xTy1M8+07G5s/oAuVRM+HgI1Z3PCMJg21piJPsrvdEGOUsv87uSmOVmE16/Xrf
Yz6h1UT85KLMGgoEvyJWW1L0vVx6+i5OMsE/IrT30do/KxFmEeN1pUvsnhXjzj4V8fLjFhouJWZ+
X39PsfbhQfPEdpTDGD4+EmOl1WZQgO3OMRn+Y/vSJkEv821XE6ZtvFiUjdwHXHuKUw5sGaBHHfep
mlPJg9ATT11oJGaXq6Fa6BM5KM2UTWMA0eMoKqMOJSbLDSXen1TCYgWEZyROiwA+Oq5AKTMqoT/5
nMN324mB6txoqwy25GKHGy6hFvLkkxtOa1wrZFqMUtqvcM4jIp4GjtbLeTB+9vv4a6ASmXOsNE7H
N7WWA1A8EPGoMYjXgbGi2cIOn1tyq0wmcqSbQldFgVlSj2O4RlDRnxfqZSiwOPMVbTMqZwttelcD
Q5su8+gBHh+mIrMlGDrWSf/4EQ5PacWySPxyiCiIanQwkiUs+1Z6Dz4Xq/9fUIRmZCudHqN21v2w
73L76i5sqQEyifkXV/0kHjR1aDdSMmKWTlduxWeuI348+HITYQ4enfKJTD8TwXnkTk17wh6USL8T
Tt5V+SNuB304/RoivYgC57hs5UnzvFAC6KFUssL8KHn4AG41hjw/4iM0P8GyUJ2tYt3L1mkXM/p5
5fVuMc6pPTOXDa2FOPrfcVriKQWHz7ldlKo4piJSMcyecOdd3xO7n3hZxkzFLdpQhrQE9ysiS2vg
3LHrMl9kdhuGprY2BvzcgaCwDnb7r1ThC+NyoKbrDqrGIz5raNhOb3Ek4IdWbv7NBDauls9b/JPH
rilSW6o5JadZRxrj7dk9cgQrBKMjqPVKlxfNoUFz0HWP729HxfM1dI0UVhgKx2oSsdPWWKWG1RST
T218ehIzHaoQvZVygtaIrsIauWgAQoyDwwEv3hc49xl9nKK9kX0UVRJyngUPzeH0sRv4WCHkwqok
kIP1j6+1giAO+jIfj3bbD9S+w16RVI07lbNiOsj+Az3whK0PMQrG1C041QNEyKwsXMq1oB6+ZNHk
Kk6MVJLx3yz65guZGQpX89cq+gW5Y63aeFprhSnVHavN07NryxL9heV1PWMajiy3Km63YkFmtvkj
OYuOpmzwvHvSPtpd1CSd6e/SBwGnmfLPeoDUv/mkcs9fGz54JS9yl62e14IKtv+uh7FH7nI3PheA
6uNYF5PvvMzDv33JtTRKtxN35m34sHOlOIxyMU7/oAMXLIsfba1u3a4p4MbAtpP6wF5CIc3Md+L7
2MvOp6GsY9Dd9T6avGOV6Xo6ALqBd9QM5exZoyK8PetJjQOrUIQk0cgnM31vjFUlVhsM8UOZo7ra
wVS8Uh0ERXkHkU0++EDRSFUeRxBL1jMan+odFUKFO+WWUEEmUBRWuXXAOhsC/Q4UCy0HnTii2vmr
4ww2+TvsAVaiuXKZ0DR+tugy666tazBQLhOrbr+7CxB/r5BmVLmAv/lTv+v/8HwYAjnkfSbCzsn5
nWdQEAdjPrk6Q7flDDs3Q3e0Ms8d72BgDS/2mCm7OO3/WB7vdF5QpZ88QClM9JOq4xQUQ9JKpf72
fabf+WxEYF2GHHl5PqAoCH0inKKtrgEZqdr1VHB+T+stjaSf/Y/lHhO5m+feSPh0ffJKSEbz+L/M
7ZRz1GRGvr4iaDJbo/WBd844XuqHB5W1LssqiuBFNn76jXI2eq6ZjIkK8A+/ezJm6VhdQE/hCvx3
N3dlPQJrY/A/6eY/gMe7GowwrASCVoiMnRu8otCZqDeAaA5/WyJoIHrhpnru/K5QtKwiJ/elgvCw
gTzYT9Lkso4by2XUc8Z9idpSfZPS9an8alp/vU3wD7fEr3X0h7QiyRKNrDNdu0C0+KFAWO3UIL5e
C02HJUXIsjPyu2WOAA0Lk5fTutQsIdMUUBqhNTro/+D+cdlbeFsIGZOBNE7n/wSCptqqSyj3Wjef
tqROXIQxTEMT83KXfHG6sDXAn2whGfbf+ulVogMgM9pnWgd49pnEERBSzbdVOKcKFvgntfXbPpaI
4PhFXDvQbMO/CRTz6ncQBceSg7eicF45kkiTwoE4Bon+oT0V/hIC7vWDnKY/zr0ejNCB1euD3QI9
e+lNqMfaZ6vXSd3ZORm0hqzJIG7YlL4E85dMviTdtacoAOMXuuTLjpxWriACYGNCAJzsAcprAmvK
HxR7pucNIxRzHgGqj6zBOzfzt8tTaN86POG1C0i8J6mIoZZJsGWgq5UewF4Flr+qIVsUfAeu2sHs
Ge2ZD83ALi9SMKOPT2XhsKE+ais9TdFL7r0ScMNDu3LpcWtSQm6w/6qOpg99qJNCvsaU7wobct/E
t76m4+kQTgcrfNeMYt3RdGuW7yqZny0te6xpuKZRjXlizz1Dafvq29jR4+RpfxrxCMaIFyTspQ4h
/RXzmg14dG6lMXjZVgRexGoeqIrNJ5drWhbaIYEWBuJNGwURTn+hBdywFeOJL3SYUF8+dkxImmax
/lTJCQXCRjrvdU+ViemTcyBARG6AcUT5YnPpnUh5JMTZVNf7Jj39zCiutF7SBaME7/sEUeRO2vbb
vjGxT4wouv8BNx9AvY1Zg8h0zAhbbEvJ0jfpBOjsssx0Hzo3ToMph/mQ2BQ/lfc5/Ag7JeEdXmy+
PHdrDdO/pQa4ERUymkhHPLzCCAqy4HhhlYLt2LtyOjBgzIDLMV4M7QhkpFUcBbWBrbaBglLUN1yq
ZPUur2vi/lRgA7ShdGYSEYbwPDk06p240tne9xWLuf7smhV8SUXs1Gu13wG3LzxrIG4bNxzV5v+D
u7a5cl4yOVkXlP0UAVCymdCJ5gM3ctzu84j+fGGwxcwcYdtY5u2YhKEMKtC7z2lzEngxxnrH6WS0
W0/Q+GqowekQtLVLsb6lOM955UTvtYSjjfJxb6o6lHIEQDE6LOl8PuHmXsnwBH/TbmW/lBfHhLti
XRu+cDy/+EcFL5nyXPmqUo5lLNLXZeZy2yJE9BSkRFw4al6Zeyv/2bImWLCPp+fMIA6DK8vzD7Ux
SaSbKr+Fw6xvjg7KlTanCCbzpzmIaKoGHQBcWPhWGc+RBMKTdfO3IRMO+xOoMI/eZWBUn2VI6XdH
GRntiK6maMoO7ZtS4PUkGAgh2JzbbMG3eSo1Mtg6KbyzVNl/tpEeodoypZzfP4chDX8UYhYeGLhX
HfIoxQIK8BnrVAyqnA0AIQ0JeCaO3cuA+jQhFlFWoQFRYmAxLXA/ECkBtpM8y8iUTT7sq29F++xi
+Q6API+i87CHKEtnRbWoYuJDoRTtMIXyLlt/Edm1azGEh35OUlKif1kXw0JQa2T6OzRYpwrmtZKR
9uMClUfC6NaxGNkEOiPKPvsSOpXzcqOX8eyvndPgsisTVRA6R4JF/G+rCta22ey9uDET0Kwaj4XM
lY/gfOx2Mw0h/LGYA9iSZ2NvRmRzDkVFfmiRL9rrkfh5rsqJ2qQ0bkOrfCfK1qgJo7vBPATS6eai
/b3ZrzkF85UhZW63087mq+ORP1faEE2LU8NMeoVOhFE5tMzcWuYOMOnGa0ZhjjjNCDBjbnJpJYU/
UrZWuvvGdZb+OrEWESxzhFvTJbnBA9Lwpw4xIjzbjw4dhQ6X/emTER4n981a9a9OtTl81w75e6WL
JoENRDvZpjPvQ8Vl71U1Y6ZMkw+Ck5dcsVZRXfpEj2ZVzjMqVdeX6vPkefFSGCUKUFoEvV1qzruH
RlSYWaLWF9sPo9RbtzbNcc1WtetxY/fDRf5MK+EDJTnAa4RoJd459wto65q2ghA1YpUaQW6oNDbB
m/hExxGJ4bfzN1vP6WgHop8M3XWWs/t1LajhXpCBCvgilZ9zYVk40Ht5b201Jqw9scHTMz0zZDWj
A47+e9dIgh+nJf52MUtlWOPbX4Rg6QtepDUzuR7RlIYxamzG05Pd12hrbDpRBI98BBfPi++Mj4oM
gJI6zAUfXkN9fjfF8K41ctpTLCqRRuLET/z9LG9AakXeur6cCK/St6rWzUIl9X2K03xhA7b1ksNL
NIjzPEtOuKhSnTUAAMqjv9rvxgwizLBDSGgzHYy79xA+eSr/97qFHabakZbN18uc2MpS4l+ixazT
yp88euvazlxnW7owYwI3ytptvsoYZzgofCSyrmsOnKDSYiEw/F9VtRapluA7dVOn+bIi0M6oHGu0
xSxpzbN9D1gVY7Wjirxg6EIYIiWpIbx3F1iw89rlluUKnKRhCEKTwvQAS9Y699VcURhmo4uyXtlv
2DboCMGHNvBsbYQQ7tI78lFJZxhlCwsR+S+J2zQRtbDKuD8xvYt00i+eckK8BVZT46X+4CMsyk3y
oyIIp0Ytln9TKRKJ12z7Rs9w4QK80AlyDK4gec0hCdXy1UwxhM3cRRP3BY5tG7s2C0WDDichRRYV
/E9E9ggog9eF84ygKaaBUxdA7xRIqQo6Hau+t0/du1SrzgHBq3dsnbxGBx6VRFgWVJzFEEgULwXW
nYhT/Rzs5pQaO2oLUcUHEHO4FQ7Ak2eTeBZTukF+79DKzNToM4k/HDaZauAQkpIUSwG4t55jevLF
HZmaVhsbkKDMySfCS4j7uDC4QUBXTgKi8+PGJyNbqdBxr1qjDEWi/dKyCQ+m+ZQRM+7zToM+FJsC
o5ZlRanUxp4GLZVQleVXRs3I0g2ADAAGJFnr8gdXbr4kP/pKNorXTBAKfMFSAfp8tYMDVtFvZT3G
kcb+r/07kZReqh5uSLH6Ys67Jef8HS7RWvEp+MZc5QEQIP+4lCQVYRAgv8VsJzAy7mz0kYeVWZyD
HgqcEEADOOZe4yRVm/D/ohbdPwBCz3oY1l6ZIKQl50GQk+lwyHtyhAibFzrbyo0yaxz+ibRbnPrJ
zr/a2aHUPR/R2VTyd0wQDyuJh67xMd56dtkXwCdW+rGTjD7pVaGCEgDhkSzkNGkVBItTFkkaxrEZ
vawb9BI0IMeDJt3wUa0op0HiwrBLLPrnZ273zPpXU9Ss12po6kwYB99fykEthdv1Z99AxQb/LdOH
nI1cqfXrIOLxB5irlARxDp/+J/LBgepI8p6mrkX4wTxlYJnbbJLJViNhHewuB5vr05M9kCfkJz22
XGalTSPPjkuE5/Hq/uDo760udq79tnObihksTJvofIoqB+DYx7blctfhi1+UbOJLoct6YgdJIepD
O53lmIEpzkLseVdC6URq6hnANu2+kjQQqujIlaaaaf4vzZocdpDxMVhv81R0wAgdXkjexpm3A5qj
zqqljHHDzdVR4obczU93ip954Oo0Bc3qT2Il9TSfMcdRxi9BZ281v3kbkV4cCByc1gj/6ls0D0Nv
9AAxc5Q3kY4gIUAlX72xWheZRmAUCnzhxRX6oimAQ9pRGOV9Rx9AJmNz4GoLA8fU5ky1c1Jhhqir
jNZOkVFtzyazOVor0dOxFOOrt7gZodOEXgqdA4IlpJpTuOZgpUH8WIjVBd5J6MZFnCHEm41TUDB3
8vocKvob0cMnbCK++IMNd9q2d+IHpzMJn9+o4yB2fJUwxgR9ALHUgcNDcsw32Mwrp2xiwPQKQEAL
UpI77lOaApetNL7Wip2DNZG6rZ27yyxxyGgL3zJ5y5BQXNMbtRsKABbA8/0Jk47ybQM8mq9cSRRl
vcrLsQW6PMSIvw+nxczgKmlIdZwt++f4qgGBQf/1rSviCKUN4Kgw48RNvNvAA5U3GfQ3OuLB+cZq
DSf6oGrlcZAS5UHWxtCT9/PAjZ3Qj2jPbCygRVZe67uKTIB/m222Ty3DXImh5EyCZToMqmnvGbgf
iaFik0AIydN8qc9ivcTxZQFetYauh7qxiawvHlZ9G70ECeQgA/7lpMGhLHTKrK5yQE2IvJetjDfU
zsu9eyA3r+FE5upf1/MY5u3h46rzfsFLJ6hSlIVpD75sDv08AiNdyrprZWfn3nNkUfqX1jlJRNXc
7SQv482OPnZBTG8jy9W48QbHsnEioT9ckwqcPa5XfKNNuNYWR1mOLDC9ZEXayS+9h3Uf9h6PW1CM
TNBv2mWdsVEds8NjqfVVmlxJtre1O6tI4/1sb/KU5bhxwCtveo7nwfJ0rDS4R0R9+mnsfsUjqa1e
AG2W7+jxeyqDCOnHClaDuAJwLpfSq+ezRThIQWU0GGK5rxDIxEUDrfJrwULx47UvQBZ2wkEjUyiG
aUxeK9CFSzMbeUfRjc6WtmiZhKaTCQLXB0XYkGidRH8myDSJAL58ppdKIMv9S3pHemjy/XI+BhDw
zDrKdO9S5ZLbWGzrpCFbhsfShLJaq7KiLAk3rvTTaYeF4/48wEEdyqQ2UTh1mqySwCMGfYwKRTuh
dnBPp9C+dYf/JYIFEQZRV8r0UQx2PeBtF2ehRvuXHoXzHFL5rlD97yF7SCSo+CO+k1WOoQeEp14O
sOM8qz97MEkf87pPaVnBOEKIhJKUMPcb2ZqXzmWSz++nM6e8W+N1ZBwJgvdOCEOTiezin/2ZhwyN
BCRIiEVmqjx+DYM+102aL7oQrACPG967l01CKbcarCrQhdPRbeiiJut1Lv5k6Gh8dvtDmid3SyW0
EGHGMHbMqm8tczOSHi+cmNmh/I3R1Kria4tuzEVROWoMN8IifBAHN0oh+nW50LjSVRxIaW0o9+vC
bOC9wGnWVQwh2jjvekzYGo2tfD5TKoxSueNgyOwgJ3KPMy/8FE2QrAbNV1KuIGTsC0RTaWDMqp+1
fIgzt5uqz6QY/2U6CEj4rkxRlc5e+mTiKllQdnYcqWFNNjflMHkli7Fpu2rqdms2fgqShDaYCasn
Qtku7aAUL0e0JjQ0JPz9UtUUcoNIjTon9lB4880j1WDOsWAoFddgHDG4Zw7E+LJjpW8qWnNpu50K
MnxrwGHHGTnnAcS9HOZfPuzmKtug7xurCWgtQZ9PcsAKGXoeD6DWTfFr24KADSJqLFklHaOSLCJW
P1tU6TxgfOCB9yiOkY/CYE/Jgkp2eOw0+/hupvtdfZaaEupG47m4jOMDu6svKsdL75i5tjBFSAbl
O/04e6uoClYdFZwZrqk233nf0zG2PSfGrfZ5b4dhPcIROcq8XoxiYne0sRoHEOUrziAPZRTBWXXZ
4yJNEZytXsRr0aQV+Z6xpjypfgCWu8rQtFCKSycja4u2wvffWTgr5WIuVXhDchGm8vUMxpV50z85
0EhxTdN32xUH5xGA6Gj0v8bRVU8Aw8tcqoa6Rjl4Arlarkdhzt1o3QeQWWv0kfmWL8ACqrEEN+Hg
9pEDPyCGfeKbA311XmzFK0wZSo3Mb9p0I1oXFVlLWeA73N0+wK5k/wiQc1wJXYh4O+4BgT+P0oDE
2zHXXxkgv7jjNg0hTee4un6iUVCqo9CAOKaR33qIP86Rw9bwvjvRwQG1WZ/sT6QY7+EDG41ehtXP
WAhAWq1WbYEq1202oSVgGNbI9Olx9bh3bjLIcUvBpw5wUabJ9+4JoBgMcbNx/CHzXa7gTmj8cjvO
hNdbgYFTlCzbyyLsc9Hsae3ai+mH/NLq6GebgXIwQj7b5ttIEv5r42HPadgzYlKguA5VqLRM1Y/l
dt8hw1XR93SrwJhK/x6JlF1PmA+HLyqmzL1fH8QfHBOCtJCz6TWZHtBmIzjQWQBy75hbuGr+bNqy
goBfjEQHMSuFslhn6oh0ITt46471uz6SVJsaKAGlrTI8Jz17ZRB7CfPl0Ou9a1l0xId3APSm/amU
KXlFlYFSzm0Id/OPjp2Bax/tEpAIzjULrVMNyeam3hMwg+Hsz4hZigj5KgZqaQve6Bvw6NzsG+9Z
hInuPdVTNBx7pWVifnjOXM2VFa0O+WNUOXWh3Wz6yJPrpgc3t395Z5ODbkAwsA94Tk7yEVwrS4iD
r8sAsOId27pCJuDgaY7L3iyQVHrjQ1b1BBdkzrSCj2RnIhOu37cgvoQYGrDFsctcyfEOt2HzC2MH
YbeP3z+i48OVuhLo2GE1ORW7ECPdwJEKX0NDKSpX7CzI3gaRnDRGzNs9gYkQRblpNmwRjCrzADhs
GqBikokM5zNdPZ5k4GK3k7HpcB8JiAZ1I/OS0xIQjLac6gmhjxfROhRCwLhsaFXmbtZEkFJ+jkDb
H9rtu5avhWwunJniaely2Oje1CVLXAxCDT042/ryEIx+ibsgIxoHB+va2OfhF4mvwfJIBFm3ZuNt
fh4k5o2FEswdmRdb3OQMx9p/1JL4V6q9SQawzJ7cas3BpzHWazyp2/ojAfzL/MWU2B9UwTI/VmhC
0gWSBINkMNvEmEszg05icL+/QpspqrzG2/TAwDksbKJ/6141MP6/GyrA87zwGM8+c7jRsCwjcsJZ
77WzTeAn9OnMFVw52exkR/GU3G7neUbaFFSLHNSp6uZQ9NxjNtYfXdkrD7P+tqGxHk86YA5hbIxS
zNMcA02mqIooVepCMVMIPPWpAkk944mRX9oCkYFiNC9ZBLkVdHccvGTMEu3nJ6QBPZz2rHsvzD9e
iWp7StBiHRt6z1KWSEkc3IehkFPlG99lKePJDtkmopzA4/3uq31+iihmTibTn2XdsDvt8bpPmrf3
TrYYyQp7Z5znW17WEM4iz/CKwf17/WPs0sd9joy/ZHjQqDYC2YadpxLigPSu9cCG/VkQaLCS84z1
R2CDdYbd65+n2fIQw9CM5LPNa1eO9IXJeUzpSH9SzG8Hik0x8OuXiyoPMZ6vzbPzDVXhBGec6ZCi
KIdXQ9ExsVFPKACZb7lNnk58IMLzv5o9GieqO6T6frAd9wYztCk0xwilsBJdBwbnaXh27tZyohsL
hrsE1F2BLjmOcN3lSmqpnqUI3k2bH5Hw2+QzKk/M3H/DLFxSrYQk+ErQaZ/h4psQTXyf9dU528cf
YDcPR3h5Yr6CotOTQEPgbncSR0ppbuajssV17gx/+Ib14o5eZQFg6Hr6B8ioMh4zujEidLm8Fpan
Trq7EiMze/KAJbl2az4sZAi54Lo+CGr3CKNDti3C+uMtN2tRYF/RwidE5wRqQ5MJsVmV3RlgYjqR
1YE+hg2klcUlc7n+BAuJQfkeFTkM+iuTaW1/qSE7RXkFqSAQmSl7hv96Q5kZ+K2w/Nyakfpg83/g
zdbINRGgtvwIfO2ejMDrrZHL5ukYGNpJ9TnpbYERa9xX/xmni5e0apocRgABIu5Dq1C2LI/MQCeO
2QvoBPm4MZ78uzlPlbzWSxVa0d9qa44Z8S76bNMQH1zo5vafdQptluiCn4Pi/xyVq2JYerF1FuEz
EyzXKSAb4/8IcBgEgv/JZeP3+d62J/eMTr1ZgAA4aZqfxtaozD/V5HAv8vecBWqSD50ciEbjuQOw
pFXs7n8dxgdy6xiRNvxGYqt3Kh9CO9gJBLiUM33cRRZqCn+Y6RQ9c+DEcjDpHAAlA2Ja82GWlUCi
V9RW4/MQWuO0tMTwuz4kl8xIyQbPyx/KJhN1Wfpo7mZ3Fyay3xNLSXA8nWayuJ42PaiR8yDc6h5e
X3dYnkp7h2AlwFynfKn3mQLX9c77w/DyNqQGgptIKTsLICo19p+q//rUmdc1N/SnOGhXyIoth35m
38MT4FjpjSvilQ6hR1MU9RG1ZqR1Ym+6eaVBQn4kAxImK35ysrGpYywb9HRecT8JjTvksMRKlAWz
H0met76NqWjjbDqTb66oqLjDBfec3m2gFMsw8jvkH4aBhINhmUIofquAVkmm0UYt1kt1Ugs5bQiZ
/j6yrDltTP2lzuDgZMKLlPTotNQdtPoX0233Y850msjgyWCX3jO28rcv01LIPWByrCRfusUwFZVG
OkY96X53iRPF67beDitcPqiC9a87YY+lFtppjW47ncjddP+HA8joDKI9fOV67YVjzNwFUcGwMXMD
js4y5FdNnJMuQp/o4oZxPqNTJ0kozLXtZgpFhPg6wBtCpQtoRY1uhsxzFPwCs1WkIGm0fk8U6NEN
jMW9yEH4YqrGAQyFkmse5+u17Ei/Op2TKMKdXlaHmLP38iS/e0raDArRmFkSfek5HRC8fYv7TLp8
FpL1jVARB0U75cAXuL4Am7rjW9wlqnw/18X8ZdWghQsjfYVhB9GtdC+SqtCPg73lmABeShsEXBfd
73/vfZcKygA4tRkDd3OGc7RJnTBHkihsTXugtoNKSLy7mqr5stAH7YJVWLXbcjX2IQElNyMAvfAr
32A+QJRQttQllYQM8GSH00RjcSqIutoczBeI7Rxtr6oxIIGlMjFVsOb68MUVuISLNKDs2DkpL03U
A4V79ELeCIn8truYVYUocr/3cN0rQAr2NSohaEpsgaVZMxNgqwA9qfoJ7QA5oNuKh+q3fOMQ/ZYn
+r4L8VESsk87oGdARIKkrXVHvHr69EM/pxzjBZFWo674WDPCIH3Pfem6Ox3/gnAw7tpoM2NTqJRb
qCGKPnbQwok961fYj6IDXKh6Z4LrQ1S0s9jBtFs0gDRxEqPjVWGg08jyLQI27h/+DR7CH5CmQn3/
74ZLODjJwPGoDjZB9gz+dyLBz/YBx4vZq0O6LwzJggd6ui9C6C1/8QoSbBahYknqJ8gM/usUtd9Z
xteovC9iXpuhOZS2imqfU4bf5bAH134sRe8VUCCnlB18+VJoaWK6BMW7H0xCr2IPNskPwD1ysuDg
lY6mhiEk5bXhhFytKrtXSGShSd6tx3ds/yw7+j5lxn2MqTEgdCGUsRMIuJJjJ+sq05M/PNAzs/Gi
FCO/jcK9aG733zYxbAzJgYaO10cNeeUWFo1nLyNppjWBIFSrRkWcAjxO6ov77HZ07J2s5QQsy6Nc
E36zz2ifrJZKuMdQ248Gs+SbowlxJ8M9uo2UWJ8prD6P4s96fNq5RvQZJVg3GBE1RDwlmUKzsjSh
IfcYlcIdBt/CeicGct9JTvSaFK+wRb4XO4K/bIvorNYKVw3NQI2vtCcQQTkfAUWjDDvGn8AJPBs8
wpf/507wnellxo6I3kSkIQrH2dhZN0eEqWx9BkuHSzHPM0ODSAQP3yTTI1j3glF/fYVzBN33B8fT
zH3ReiA5zdug/ja5oVixVEO8Wbzsmq365shsQyieJahlgsKpFeNIioBEhDTNpyTPPf2QfUc7m/V5
kzkbgXPMeaC7RvgXes73bCwurubRMcAqCNx1LuVd2tZwnHjPed9CpESfqBEkdGDZxmCuasZANWUq
7Rj+4zjRsDCtR3gFjrkmF4Vks6Lln3I225Zaq7n00GtRWGTBmjst0WlOOvg979CZBufba99xxv+8
FYyQb90aMf2G6Q+Hefc/U4GymVavX2ipwdI5xruydRysePlYdzMbe4vJ1l4TQrECoXGePZ3t/lZW
zBfpWiPs1wAMKCN64CFAcsXc+Uom71/70P+ovtRYGXW6SHvJxAWehGqQbeHjV52MZyNiSUuCU060
g1u8ia43ML0tYy8nk77EspAGo0yyqdgs2e7UwC4AxXcXv+mqWv8X90P8Hv2AlvGyKqTtSSR+4W4j
ZhcOh+gvZZQ09NPuVTW8ozRuYmDfCCw2P496O5aTwJb/iOv5/I9YLiIjOjJVqoi3POSXYoeaNoOp
1Q89Xu2XnTRMZWVZS+Qn2TK4mepdz641xSfgsOBBhxUy6oA2ZZkq8QqyeI6vo4RaVtoYVEZO2vod
Ve5vMKOiVMw6ziCQY/jSwmzbpgbNCZpbVrrrX7eDvvga5CVx1Y8r9sEGFN7pHUGO7zYPaYkqEJ+Z
6nAP/fzZzIljZvl3vs2YtFdk54bPXrxd86hTB2gPDkusZBWxfG+Og3yapaulNzeriyWWYNyM1+CM
SF5dpXWOhzvYaUcmY4+tSvq9c9lUqbE3SL9kRlscUB0i5hqhOq/7HhHURrFYVoUWMpiRg70F7qKI
02L4Nt4/HjjFFB9Ji5RdJqHepRJdQTI+zC5GpGbOgYK8/S2dqztT9QC7y5PX7cVtOstLa6T4YQJ+
/bpEVlCaZ1ZtEg79H7+/6YgIrdScqJcg5H5n6dEvm6qIRXTpXA+yNUhxo+yyC30zL7DUKH2iJiv0
qlPzOQNF6zS9ft863KkLTDtjadcEckd6XufAbAEVTpspHDiQwdl17z8lCfh7huJ0vNpGlX9j1XcD
qGqzqOZMbC0T6xU/4eBrrUm0dryHt3nl9Q8pDZk+AiN0NObugxueDlBUWmGn2Co1T+OrKYrUt0fM
tVBPoFbGhKTwp49Kl4fCLUauQzYlAZP3gBDv24rH/AVCBSRm8/V5TSkTQmcNsm4OZ32cm4cwBQ3N
Une/LX3T30glpqW6PS4C9TKQ3SWLwaOnSpH9feFgxBw4kTTSLWrgrt2LeK1orGFYrv+gq1NWVGqn
7LcPtaOH8yyL69ig8V4RIxKshb2D2KITp82ejIBMcpjziuIey2R1lgJJMm1BSFxqcniWG+fY/TGO
3+cZne2ILCSsK7s0DNC7UvQiAIxi8Vyqn+2hEyxLjCHxX+JWc1rZk7vCLc4gl8HSqrrM7A4pz5jb
+6dQOIN0AM61aReXzJwDmrOElMnS7og/luGuqpVKPwVFHD32uEyz7oGSaQZZT3NzzB4jLmHIOf4r
gHpcHwx8XN/J1PVlXdrXWN5x2lUC/WUpKxmschZD18X8UdgigAw3g//aVnFLaKZp3yrlPxLslh/G
hdrAarmpgzaJwhrtLgBNYJHKCzhNfxGySdH8YtH7Fg8k6gRYgIf4DFZ0B5/iZd90grNDBDCk7S7f
k8kqZZq0AkTmErCSfpphJ5H6AObcuxh+LKh5C/09OEvm05gnLpN4cPkecXH46COnNgEBL/ifFqe0
WsxxbGQzjKdJfpV6aCs4JO2urbhZo7oTG4V3N/518bBXN5FtR57k9ri3IRJWX4fPjGsxvkLqOPyj
B6VW2VaoB+bdnhZprWuMcOjyFB3dBf7p6XzPQ5kdgrrsgN9MLpNKS9SWwAQE9qMoxrcjJ2ZhiZbH
tias9JaZkAws0g9cGFzuHF6CqcuCk9fw/w/vk+oWuk610CCItUzBzfUUyHYh6Dh4QHyUW9uGoRXd
cvFzZb0kirNUD2XXQRll8q87vsA3gBWSefDPzWEV4HiOSk6zElYOkHPKU42OdWs+5EEXWbaNqb4l
EcrmDVZutg19XFHDEvL2Q9BKgKnTtOYEi9PKeZyHtJDRtK82W1Svf9gQ6Uo4LCDD/GSLpjSHIWrM
vhu4v29z3wlDke2tYHj/xH/uC5SJic16K9AR+32xtZPyrl5AHRMCLPeA+Woh9qKb+fxHwXdulGDR
M5GoJ2scqPHh1pjZsDXTA9pp9/u2xDaDa1bIMerUns70spjbJTa5FbJt+VE+DVKgvOx52J/Paunz
39YySNjdzBnJegC2FIBFB4G2YD9HYBvmSp5Az2RPzcPmEqeXAtmfTvWXiBXquEEC2YqutHm4Dt0L
A4oN3izYIIHFrBKOT3mgOYTJlNe/7tcAlJqb2Yh+VUmqalc1s09Vr0pQBCBEk3unAa5FCverA4zY
vYQARsnA8Lf/kXGnl4DW3m6qX1r8TqYM6l7yBqOkGjrWu4KBNgM7EBXy1vIlrLIQ2IT1tF7vToDI
t/US9wCT1ISjVYnaVxsWwmG0hxKKTMQYLDWwYZDP/eXwVvQJtjuhqPvirailGGCfY80O/99fD4ue
dxAKwot9AQgbail3IDqRX0KVx9S1WeWraMkrvASbI5up/HkPcoLcckA26vHdDFseDaRk/Q61IZgC
vSXXpPILf1+s9phj/zpPlIB47BiqLC6LgDbRk51PCGSbnw1j4OJjlh/pzWF3dhQGYjEn+kaS9Sif
t5XsBhzEeKUvQayAFqzylAPrEL/+lbr0BOnQnp1ipNAaRBzqkmLerX6GRfHPULSFQPk+Z6duB9AN
w45J6UXJ4IhHmGY5+6ZCI80Tn902KKQblsXZRAT7zPpPbGebwWo1IOCAV/RWGSRo8NOghq3mMIsv
KPK6ZLbRNNzN3WxRSfu8MFMTE9jgdwX25hPBRp4i699/i1jvVfim5e4Q91hAti4AVCSs8HyK+fys
XBdHl1mh1KNBfJNPzIXvAIPeyLkjJzTdvqi82vfqVPO2eOuLx5Pm8pjcHQAMjUfI9CJVP9z1TzGS
O1ZuHU3ILXoZDwPyXuWVQS/ylWN3AILhbzn3i0NEKq0jTBlwuoMmO4gCTNjKe0IApPu6blkhdiju
+LgxxTVOGY1Vx+ubvomliupKs9BYMdVEh6gNNVeeCeG+71vCBXNmFQ3u8RPwd+WVbnfExnIZMzuG
Kyblke8iK9KRkXH/qZtmN8NlichltnWfWPl6knedPSQ3Z9A8PhH54MAG1RGFQaFKFGXBq7qj4dPu
C2u3ZIm3bUs+l/EPkJhtPlzQJn4tEFxw4jvbML1SfZGZzFtCzE7glYS8XVlAkizZT/eVASYp0JvK
eI4MyLtlqQk+G0vSzDkAbfmzs+rMsPGlCasPPzyNP8jMoqN3aZgDwsP8+RbyGU7t73uVte0/3ISS
26Mm29A9drAo2/mILZWGxJmyKeQAqhIy2Fg3tOh7G2t/nCqis846RIyaoku/zLQXp922c1dUbAHe
BT49xfM7JwzWyalqOtGS3O3UWPg0NU1P+K8W0kzH4dRj4LSMXURPRUvN20utwiz9rWPWGvvIh6pp
4zq5gZxF85nvoio/x8LnjpRfu1sBVSOHa4fuTqnztFSesX+zDZWkPELmXxSo0qBZeaEmXLtITJ/a
qGXxQp8OF4thDlsRYZq31nUvr3+HTlzRcYPg2GgsQoTf9Q+hetlDmPbjshaS0QMBZup8yZT6rSYW
YwT9dpmxKmsAPb4MTHKwzE20fhhPnU0WojSyFc9SBe4kFFvx7A2BE5zXfJf1QeAuMW2DUa+l9a80
SK7p9UYhj/8ZbrcW9WE2Jbqyam6jqlr7FYEshZ+lYZrSITyrLVke2x3M0lWFQ3E68FYYNNK7kqEx
Afz8OmUcHnTQ5nlalshP07b1IVFRpw2g54AXTOB9TH1GRxhESsldnMJ2gtV+zupYFYXydU41VPR2
21MVsdvZw1vw47GJ35Scbg/XRea9yEhMu7QxwoD8RRoL1vjUuosYyF8OknCK5URDfA7TWZpSh1K8
KS7Y+850jOLMzkQ8Lxt+TXEVgt9RLiQ+H/xqF7XH3U2zSE7d7akejQFbsL6O+RbJXRhSA9fQcRoQ
52/Xh9zBoARz11y2nbYVw3MNQc/UMtCqJxH7X+suKeLDf3JRDTqrvePWN0Pn8BKBweMhDlv/1+tn
vcMx+RpaSNlLWsK4LEIbl0srEU86PL6eXEW/fdRduGc54vOnURkTj/Rxcfi/UM+OuvO5SX1JHTfk
KSJBVM0TZYBqhAdHlbn4aTWTmQUXpF4CReuBTIvWy/SczH9fuqR9GIHIdnrTdquWHsZ+vG6ZkiiV
u2gFldtyzGrd1ZoDqU3p8uFF/AaP7Ot0SzQI4hgAkc7srksB9+dHOd8Q0gYXZZCIZZzxb1P/tOXR
oe/g0n8BhqYi1Oeunwx6EV8DSnLm27alJmn5z+j+AqgJiDf1sZjTVjmMgF8fJxTpkkAjxO1K28Ve
8Y1kLFbUNzJ6Ro9hAPqPAsruLnV5ntU6TvSoRO6mcpthRt60z2+mN8QXzZVt+INBgvrr1haOLrSO
CqdTyXPi7vPnshPHrMYv4O7mTp9u9Y8WbGCPh0O4AXOYSzNRbANcO7mEnNLXfMMk6zAn4MTI9cE4
l5GOlPr8siKh+nncSFUkqE4GXq6jCVOf+SFfT8715Jy6Ig4VxDD3ffPRfUY5/rmGirhZNIc0Vw+g
xSQEKT4/+uoAHMbf/mQoC3zS58a4d4sT3PLs+4nAumJlhNtG4Cy+/33FRM7YlADezK6yfJz5UU2w
+OJwu9iN7dANyxxinUiXK0faMQpwXJIszihMsoSIICtSGCh+75Nvx8yLHjfsQk3CVyBlYty6Rwnb
9oBukNzSwLTeHNwJswVshsO8g06412TduLyZWB0hvjLRMxibltNrdnACqkNhUrgeMrflDMglKKaU
VPXl8utCldWri/psQw8POVA8Yo9al3fXj3CbJTRQV4X0+w61DGf6DDdBmYGACTWEN7LXo9/EAQ+o
Zl1QRW1GxpBUImTpwF7oBeBXXDqN2/EfH3ThXz6EVjMKzNvKPq6YGoRmdm9zR75X5dGZXk9/Iu2o
yZdJPhPyA35/P6kIm0uu0H3u0zpneJKKmo1ASryBjygufIiMASWF6gWJ+fqX0XyyuFR5mf6GhIt+
aVhJvZnRIB1BWPf2ZuFFoG6oheDC6sC3Yufio2PopzGfPNFP6r7GQFrUnoTvaRGK/OMsGtctvVZu
OMdT712+Zbv29RyR9LFS3zepkN+aEvBStPdKutsYGkhtwyMC6jyir3qwgM8B7dSBwuTagYajrP1c
rYCJTMs27WRFuQWyA69n5M39vRRkTmTcPtD2OHOirRHaHmGmCYJziWeUCpAHB/QrziHXYUlrh/O+
DAKAAt5ZGlMIMQp9QbbLjJ6XWy1AVTXqeW7yiSjgdrH3biL65AgVItIBH+Ele9UJPAjm6SQRW6rs
WE/Wu4AWapHPBcoOGG5T8h/tityQ0UrZYAg0IUxI8c3SHcUbSIB3Q1i338hAaaYwgZK5JMCGIVKd
2hfutHSumUFR3ksLUgMXVFUlva6PM6ou8JZNQj8xehc0BE2ND0yppDVjJwrXi2x6eDYU1uqwWACg
LHD9sYkwxECyNXCmlE402b0RRh6F4Q7VXTgQaaQdBMd/qxgQbhQmKOwgYezaFsbgggu7vlRhtsbc
y+aXJTyIgbpfKdSlG6i5TCdgg31Yp33KMXkTs7Mmk+vgOgb595kv6RM1ooTcfYJW6XtkysaPYcNv
SFEYC51NpJKK7/pdbvbnsid+3qXNJQtsVSX02jGYoV2qx7LekpK1Rpv3W9bgbpH3NKDYehTkwIzL
fXO7+fSRFq41a2TsTfS1LN6z3FPXo8+/jPxy5zWR2vqlcsKfwRkedNRnn89PuQJbZPIvSGD6ZChH
3ucOt6sOM095WkNyUEqvEz7B/fxivW9rCvTdAUwLy9bVKz1Dud3uC4ZCmYkkJ5BD5KZnTGwykdiy
yqCD8Sax1hFGlX3er2e1LM10MnsuAK03alhAv26KBtxP0HpFhM6QsyfXPiE26EsXEhw+HS/byfFT
e+w2wLbWU6xbpZ86dXy9oEKAUUtDoze9MeTo+Gs2VagUP4hk87GK6rkUPJqNxL6tYRoVBIrRxk/0
7wR1xIHe5boyQ5ryEdRYdVF6F5nGNuS+8h84gKxqajsSqSCSHXn2Y4BSA5E9zt+d7bmXP9stOkNA
xXq1eMVEg8oVIxejwppFQPfXRmjIaUfCx6L4IDOA8CRltRfa5f3BgoJz7IOhtMOD/QwAFUWc9nvR
CoMfjsMXpeioRtMQjb3NrGnMq6AoY6C1Gb1N5ypKxnit3RC64w4Q0bOsOD1I0QFhiior09mbMkG6
OznVmvKbvrxIZasCb5F2VxhePWH+wWV1BSzLBW8ytJgm2t2eQ2IM3+sSAbA5oKZB6ROTnbTJkzS3
20Vrn5oI//G/pIQkM1JkCgCo/if7OxnxooDecf7GUhAVSWBPq0vnB9y+91ADZUNnpNERwfwsL+YA
sIhIp82RZ3ebWo496GbRx7nZkOWkWGE03aWdmJ0JMx//myYcRL6ENE125Pw++0kcMZQMSZZhN1xC
s9GGVpPCqi5CYE6zzIQ9KqknS04LOxShsDJiMgD5mbLfaln+bNRvwheDUz5N1a7P/P4OPqT7hbFa
E3qYSe9r2m8yF/VyJ+TkZ9lIzeUQjhqJbc2hp+pltoFVxo5dl77wdxOfD5ztDMx0j8V0H3tC1u0S
ecBZtxbl/G1FkU3NlGNFRLLnHL3oOYTAHVTqMGlG1nB0leq945px4Z7HbPiIVEOWDakgWJQ0Mp1j
f4AlLGr11Ugz0i4MHw6OwJvEt564aDaxc9vJGY2oVLyfk4K0WAHO3WJO6K8dW+XeqrdD4mLXE/bC
FEnhFehGjonR7DbLeSzNgl31FCztMw0BcPI4kOCfptE0Jdrhqoihw9Slx8zc7hbvxT7iNy2o38h6
/WreX0cGJzCyjCmk/QhLawCoxC1FcwvetJordys+KD23TTmdGNCfvCfnqat78UV/i9woRpt2l5/J
eptl6qm3ibzwy4JZ1jUoBDyqlZy2qXBaju8+iokjcw2m/foGXAIGwHW71d6YbmWNlTMHsooTT2CY
+LABRlCrMqR3/RS/6ERtAR/saLUL/jXX8nULWf1Ub8OLAeV4KMqmwc1AP5aCqxhxEZKdcrn20LKw
KwlyF1Ej2lfO1XR8QF2KrP//cZV+48VRyt+HyVH1YiRompXtMSoWkBWKFawKlBltRYGY17SKlqka
idaSM1reotU5h2gkALQ4A9uq2ZqgD2mg+1xP2VZ9zfd0APeiiHFjxd/Z6eOy3QSSqD1YaunpYuL9
AMEGx3y0/OmeHtogNxWPAZdpcPbDEqlNxer5AXacp+Dcxc66jkVfqSdO9aZFPGjqC7CToq6jnrNk
IjxlWSKQ/YsFZUIFI1UZm/5LxUv8l1l9I1VVlKrOQgvthScA31xn4jwrlWa5iqZ/lwA0JHhuL6BW
NXjrgVcMAuNmhp21UAlCIHp2YA6AhbA9JbaMAlmw3MxUqN7n0ECHSc/Atf7AzfAsORQIC9ISPOK9
z2usV9x1gOTvmg72iVKXPCkl5U2qcu0mVbsosEbLycqINIK3Ot7DAwnXkuapUuMTlTA4GXGFL2qm
R6iJkfxQ8S37iDKTOFr1xu3WgHPba03apVjVN8qfZ/sSw5W2DNx9NIuRLPcfMZFGNhltbt4EloIW
gVq9n5SiQlC9uKAvAFALdSvko3xi0vGXaeY5aUNSZWbfk6ZfbsfY2gHEagUiM7JUDJx+EAb03SkJ
Ms1opf0sQ1MwJ5YjJnWOWmUVMXU/lunH6Z7dJMZhzrj7mBaHYECzYdR2wAv4rG/kYCCR1hMXSR53
3OFye5QsEL+zfhVVsZL8BXPLBGOXYt75pfNrKGkwiNAOW2x310uyuDvUf1pkdIuMo3DxS5AReWjz
u9l9b2r8O6bnx1rjNqc21CKAa7XhOibsQO49Ou6I456IPeCvo7S7OlvDrTv/7Q4mhqxzrP2GIq21
faArUeL1fC6PSn5Bgbnu+BkOV4U36QMRRlKhUM1/Pv/7nUokW2QK74fhdMlhhH+BOM7svGG258hg
yMQJa0czBodCh+etc1rP6Kdk2qc+yquvuBBXl1SK2V5SaVe4754zqWuGQ+5Izz7p0RoUsOpmiiWV
QEIVjkjHcAknchAJxnvPXhPzHRRHb9UWw0t4EQXm/eWZL/+r2TgWKq/E7Go+m2N0zv5ECehOgfVF
3KcOTGxJGcVI6en8IjyIlbwevCnK1MLRE4ynzQ0bDhf+IwEv3OZSXoNatmZvLFtI7oxXXE+BxqyN
A62m4oLOvfxfHNfSV1672uOjx4D5pNkCGSwpoAm9mVFMuy6QdQ3VXlWcJs08E/yO3D4XGPRPN7a4
D6tpjhRq+eStdrFp3QjwyJ8Wy9xPw1Jo11mo0uxKb1qxHVfMEKhxb7jtM+LYLc365Yr3wOUQuw6Q
AbRcfWdHvDm1hIYltaQUedqIfTaWhJBMReb3Beb3ox5LtyfRXvip8gYXdz8nzMhVe5BdiN9GbWSp
kRSQ4M2Gjk3Z1bI7v+HF0N5deMqgjGADSOP7gtVPllXiMCIZC3UCOhAeVVlokU3KcDoPmhuh/+Tq
mSRoZm/LtMeZTlEV4exWBKElvD3HpPQC0cuCHeECr+s2QG+DyJf9+vB63Mb+asr1+xHCUgOAY/x8
8Mz61rwYV0gwyOe2SDMgJOeZbbT6PC8pCoy/34TiZhFvQDyCQif+qbhdQ/9MEyrXLGLCFWoG+QdK
tNhxQhNrOVeln1r4x0ThGOTpjLzVEYA7POF+6u8N/FNW8uLh7C9vGV1m050e9zMXfK3VF6drNEfS
t4ueRImU5lIReCyk0BcmrAe1L4PCiKXa7RBOPdv0UifIY6I+yW67ru0mATRhCt2l/2Jw6qyJT9be
padw3OpwSvMJc0rifVrrZEri1mGAISBoR8ZHTD1HrJ3R3xnSIw7kcEqs204PDvqgshPbzP4HvCLG
u7X09HPxD5SHXdwaoyrzl7xUo/eDFeZnxN3STWUsBzHFEDuGk/dYwaefXCoXwstqSD/+Bt+scLFz
rbf+caQELWTkdIs9Q9xe1xJYNNaEuO88JbYcTX3C9VfOxUsnRd5W4OJRumlcrmUbpSdfDgKfNJdx
mcfJ4YEKzSIa0afNCY8kcCoLVaJFodmK8shAbQ83/zpDeg4YIO+R5xwipGVn4VSdyqfXAnBEs9vz
0Acf5zitnVz6hZ40NxU7zKHbkP9PyKrOXWMm87+fh07n1/bHQgH9SqhVwkv8zLo+sy9XNS7YAXkC
5DzGr35A+NiGjsRL+bFdqNoBB94Iv5R2R+/5Ws5VOBS7zit7TsevMkLky4O7XaH0oFpWq8UOiM0H
A3nCSvZSE9Cydk9GJZoaxE+soJ4Uiwq6h0WV5qvj4Vbv1zLgnf+ogxW2IVFNDhmEaKvt8aG5uN9K
KgKWrn9J7s4Fj4921kGYJx3cimbrazAWYB8cR7132ncpUGUzZG9+WkxLVwHVYWUdKyOjbqlR3Mf7
MVv94m1fhc3UYnxRH/0s/rOVSOGIb5SE4tDUkyLm159u7r7zvyxK3J1FXctS7YBkO2kGFZMvgMpA
FMvd7v06fEmlFn0x4OrYvefmrFoVOvZISvdXx7l15cn9ZjdCwraHArH47ceaklUAEDNmoeQW9T1y
K3FpHVJjaZgiJpgHsdJjLLCRm7e5ICa7AKazTykDSLanyXaiihamlcEr8WRaUb9h9VgtprjcDqMk
0uQSnilOl+uHB/EGWv3isFFXW2Q3hhjSe48o4RBYUI8mylGdhYF9JYJPB5Z90tHug9rlq1vnonzq
wRAWt3gBvim8k0XswvL3y5mmNUekEgrSh4iYLdGLE3gfAfRbhUheDU6WK2gMMmugkGavagJPGMAy
5nxLE+yWLztKEyBXuf47T+9/33uZORp89BESlLlffpKyPnnXWa8yTrXnx1LCwNUgmv9YkULDH7sH
yvuNtmljtls5S1vBuaAnsz4T3F1VpfAFO+5MhEbB7v77ZkAmgU9dPoTBp3mIkI05s+wisWyemyTV
LDP2d7i3zYuazAkI+ac8tvfulU4ruNsh4l4A15XmvUNTskggf+2HZ5p1iZKu8dkjJtXuYDzHNCIq
g10velVHuDNEw6SWVjCIt6D4GPJvPGswmOvDd3cbO83qz4JB6hPSvwY2eq/H0yYAVp7LFzJ0o0wk
U6Y9W6tapMYL2HA/UvQMZ01o8i96I+OuSdS9or7ubdYNjkUJkoNHK20r/3WRnNCWH7uJljSvlfIQ
hAdesyajtAgkq/i9t2IBALEkOvKwXL2N8jrDu7dHXhcNhKHheh1mENzHxSJnbpYLOo/mi4Ig+84e
KqcFRyFJDDvr9FJnKp8ISmrigZ1NhbsMqQP9ps6iWTN0DywxL7KSEYIyAos1hMWClXpDJnd+KvhS
hVZICtTbajC7lEBKTB3d7kSA6vxLxaDZCI7cCzuPcpAG0/mEeCgw4ejki08KBzm5l27GfNFhGXpV
23FY2xYGyFZxgBRy4lV9u6j84frGiVD3HWdfU3Imv43nYdz8yZneYFwbW0LAq+d/eGInf0IQDm8X
BN58yA8bHC1Ul4bEeeEaPmkeTM9v/iZATSS/mmQJLxB39f8qZ4ICksQQTsjx26pvuuXf7Kc9G7qk
ye5ZfjLXrXeWq1aB7qNVnUKQs4NnN2eqCemdLsOpzZLiQpS3bjyhT1Plk3GJHB8TA2NsM8xtl2uQ
mWS/0ku1Q6h4UHMKcmK+8AopNoFzcXptfBT4PIodXHfU7DYYF443prH7YJ/QNwVwFjqIiN4PduzB
WT/JTAZqrJSN3yts+HZFSICyoZmbYOxDQ9zADTQ6BjqUjLVDt4oY7xfiwaYjOnAPvSJYsr75uS/M
mo+tJ4eKYNfjbtLUPpKw/hIlF0SX7tX1mMas9413aW3M4DaCO0hInXjg4vFnfl5NEdBe4oqWzwDH
TTYYINE4mrv8h0MdzSKAFJ3UXA8/khN6tnBueOOTLCov2A0TCYAgHSjm5Px7fuYztWH4+ytgsIMp
TKxdjeXPvpuD+J62+K35cXxnCW6MYxSjsdiqnV5SNxUBK/LmBE95phfGFiL/BIqOXZOSc74WmFwu
rfMwJ6OBwIsBxbYzbN84ZOfExpu1vIQZDqfLuU3P7LzqkGWjhT0Csi8+lTQdi6PxjGfEzD+vhhhj
U2GhVjDpIm7SAZj0bsL0/5eXv/vHAoRyCweQN8aSj6jSjMFlLcp6taXjcy6F921V/H5WfZfxfSPo
CtfgoPEi1RoFz421Vx408EY9+5Uw4hcX5yh1xfyoc5X7WfypqhQzy1UfT6kX8W5LYS/sGjAGJeOi
sQ1gRmgdDCEmpMMGOsx0jAZULV905VZ5BXMN8KucjFgG7Q/8+BGPncAxd6FNEPXqws81YsQgOkn2
xJhjugDU0mEn7g2L4mIXydG5dXy4entf4Z+udLhqOtsZLZbwLAFIbnYbsTG4duBVeO/IUcS6STub
yiTGietWcVlYnttV3/KonkMXnbWt0U7ikzgJZvKA8KafqdJiaHYhSnhq0hKMP/ze6U/4/fyH7kJZ
nJlhk+LNyKWev1IawMPgavsSHq+9JpTw71uHHqAB4R/HWPx9C5aoI+0ncE0qqU6hv3OQrctEjhVz
MFJKGjlLOtaB1BGr6HtmDPvJ0DhAEjX/3b/j+QiAbEsqqz/HwjyOrLZXYAeLw4eYYAmyFViA7kUu
F4Az/ZhdanNcUswrraSJiNuj7BN9rivUX7iaPrvAgtokQ2sFkg/7Q1i6P8Gp/jFXznCMdrAQ6D/8
mjHjtBPIvQbLF15wgTYBWDQJDnHGaqb3cQyZKzbgxFsAxsdU9m7p/GeOLp7j5kCv37c1sUbjh64g
qO8EZvzRrk5cyiznBTNC5BC/bWC/UmAoYG9CwvMKuMg0wR/3dLSzErJsOKN42qFyYEVtNWdL8EmS
vVGGz5BKbVpbon0m6l26+iMH6zcqQyGdQmWSPuQ50LrvlysgaXUqZmBYdNhQGyTV3EqhJGjNSblp
AT3M7zQdyq1mS95+tYJPVtp/4KZOxtclxG89fdNcA2e8lBOH0jKLYff9PrgSUKrXOCMTnercpihh
yu9U1cwa7/rmT+TWqDnRZzo4MhCj2MqbsgBht2OEDyUwerH6qGizL9KO7bgse9XdVSBzRLIwGjGY
aLkK1ekWl4WC56lR5wq+gQzIb8P6IhOyx+O7+FKNY+5nWwJstI/ixBC52wKLYBL+vvGKSxZN3QE6
QnnzHPjuUt2uMO+fcF3PR99lNF1zUwS379fBNj79o7HWekreYLGILZb5l9tWnDKkD9H3yAkScKe0
MVLzsLtdfuUhJ/OibJcKhFYDhdjxMqMKC7NrFAzsKEUEBGalF4T5DQ2w3T2WTBDSx53zGu0azhvM
VE6NLevcP/NgJD21jGUyIU6daZYAXg4/TGIgkPmBK4TEvzHBRJXR+n6tcko2vRM0aiKvvMbJPtqk
pKpBnVX+fwOrZKZClePJQ0KcLIiQopMJtesCPs5haUdrvvIMuNVpE+elqnE8Bv3VUIailvV5B7Rq
SIQfHTf0GRJbMUFJODCopvm+uxqqbcxhWAB5i4i6Wlucb7iTMBS63uZD9CM96Kz7vgc+a9LkRCfM
kr5G2Rn8QXsLc5aXZX0kKYcU+8Hb8Di7gV/7Bj27lZgDt1hEFAUzkUnBNqiqk6IB1ZbaLsuJUkeH
0CLXVaq8yCEDikEDVOetakS/+k1v5eNKLK2Ce+9677QlXt6jGL5bPizflZlfsUE+y7q/YG3qZjSf
aN79iN7CTmtix1a8DxUGiZWxGZBIRkTP0dTdBw8OIxcANo1J8eJGRJK/bsgN/BprI4fWsRkZ7FuD
xdNyUZO+/8XlLRu5BUNGbitVZ0kKe1G+sGTShB1wF8iyuk3LG0Z9PB4OKGGz/oShBmwxvkjug5cG
3qxPiwsjJdDF+wbxvr/VVQjolgAdI6vfmg75GFGSC7NhN6IjN4AlCNGwksrvSfx7l0xQlPO9swAI
t0PwhzTNhFQ0isTLTpwYcYyHnuCXPtltVQW5PGRSeQo+7DcRSZie7bi6zHEuV4odh0ZBqAWdIFxW
n1SNquB7Sdis1fcmdrkRSQf0W75WcjXw/kTV5Yb7AImMmXcm67cVMV8YH4EJ3MSTedxhB5E8EjJ9
q481SUtdq7oXiFowA47OF+yAoPuxTe5JojOfbVm7ITQVOZ7232AipvcemGZGsVsjzv9/W1V3UzuC
Q0QyDQ9ceEFHuDDjRZIIF/qG07vR/9jkiuafBodmvq34Kc6cCwjZNZhg9l/PY9TPJ3M0/zx+LR0/
oI8RljK+PioCg+NdaTgUVmwSfp4IJ64F6AnaA9j1EfD/Ss44dNV68yHGpZZ/gMpByrEdcRm9oE0g
bUjRann58p2P+UGxKYbRkaV6fmfZUyFdv565FWMtymrlaEHGbXZX857UfYbke+E8uirTYZXWL/oZ
SErLMA1hMPn51KfvZwJxdrvVRBJTLx1EqmbPTc8JpaXh1CKMFqfqnSCJP+KreeWiHvrzZPXX52j9
eipY7F8iHbC588eNPXRA5aP0A13UjKzEadZSIjhcPy8vN+Uv0+b5Gg8hguguKS0wbGFdCRhRr9pM
51fqAhHvGKRL5vKYNzyPDH7MsowMz1NSQUSA1obvKLnQLFJDRmN48XFleJSSXgT8dJK7p9AwXoUh
WpOLtAvEKzT23lKm4UiLOu8QlyaarZe6lEUpUIcogaUkx5UE/9pi27W/HHnfBj3n+0nVUKBzwtcs
ZSZtFzKg68FDcfwjEUtPNlZMIv0X8J2JPwSA1+0cXEyMtQJ7Slnmr4h2zi8qZIh5OrKAWMCxe+XY
+uKC3N8dwGCk7bG76/FAP7i8jBCE4jaHPP0Up+4syWu9Fym37owoaEeUwsi5kmUZAQzU+FH1ezVZ
SJqxkKNrH1dxsO0q+3MXCOH1vPL9jmv7w/p6/1mYl9sfkujztJ7FM13TO7oQEhv0YSY8EcVYhlnd
qgNWL1ZTBeItuaBvlmXqE+LvpBWDL04l1yYbajtKz2ulbFaqbCsWx1Wzf3/65oD1DZc7AWq1JliL
oFzI9CwDmWswfLqJsYwg/bSBExyl92XBOX4BXoGJqxchXSeX7P+5KhlQBHjhcL8Yh6CDu+Rpd7vJ
zC9j0DLcCDvsH8Zmb4mfsQLK/OdNQ2Qjoj1ShFFEpDjwOpkX6mDNyBEPqb7IQgu5keGEsWfmsUQS
whbSL5PNdzT2Hc2dSSlL/yhWlaZNdN77YAxifcHO6z6zqxGsMSDwTBi5+v5qGYHw+IyZ88fZeT0E
vrozXEW1JHNIHqdT0aHWoFXIn5Hnat7ZfWNtRSWOWr3CgZkytPcoaWRMDIcQVNusDwSvf74838Ba
1hfAA39UbxjEtPAsekU8TX3dJzuntr1OXxS+eLEpZvjGsknDb17MMt0neznUiiKaha9nSCjQSnXh
6SM8Qe9t3ro/C59Hp713CrZUbF20EjIv/t6F8xRAKDWdsr+i9ElGqg2C4qxAFdl+yQbgw9aQSGFG
iHqpU/p5Gp3cjuu+N9E0sO12p5wqY5DB0OvPT/05P6ppggeIDabO/wrljYy6VzH7zqDDrCM5DUkR
nyXz0/A7Wvqdyxi5tjpkOfcUiU8ntRPibx5lruWL00hgASX9PJrnSpYCjNy0d06OsEXTtFYHM1W8
fVAvot/x3/sqIPTVoognkK3RME5c5BbKIlfhgm/xm6QSfm7MeiF8fO4d8I5/AVGO8FoCzNVfAosL
FyMtePGHJUjDBAtq9y2VBmCfubJcnqws65LqdNlsAH1+b/KT7SrLpsZwCgL+MLZpDpjjxfSxsGBI
KxSxUKg49CuS5seTbB9FiaAdBdgIn98RJG8MQRFdNNAXWkhb/n9sLndpCY5RJqTmTpEMpFmmL+cu
mMLRy2Oe0MOt8CKFE/ihEj1EdbZN6EzYj/hJHO37uK2nuKmsAAFZjJH04PpEJBmJN0e84iPqbpC3
N41sgs1wRTuYq9cUEsqcQ3It2E9Lo+Wow4fWPRYBF3mWin/Tn4Dh4pQHIM11ukD45+p36ALdDOVb
16Gor4ItCVnZ5blNbKjc69BYl0yDP8LpTwUBvxpEsuISVerLSz1qqH2kEgQ1Xd8CXXQLarc439uy
ZTEL8ygdMyUpsPxjp/ZxWpnNddwGBJnw0y0UpVG77yBw0rCvrex2VJYwZewIxsEotnfebe9djmI7
kD9eAgUO1lAuKg1CBCdTv8n4RICOwK8zYxhwBm1HimW6eQuir3Ibhtq6kvu2KKScZ3OcehM+Ckxt
tR/QR2fvU16iUmRVmrDXiXfEpnMEdr8Gso81F+sCBwhKfI5Sfbi5eXtsxlBkioX0JT40aizFqYMj
zeEou3+qIT4XxKXJXFIFopYwtsWgV5Mj9i10nDL4eJKt0Lb4iWfqsJfx7WTWNR8QeKUWnpl2VO3O
5/Xw4X+/AHmPMxeX9qZHoR5fkgwitztHIUPuvXdQPE/4XKccK5/P2XBZmJEtGTUXIOiC0gkNyxMC
+iXvtdSCmtoe2FteV0VHNw8vvM9zzTF4FXO+sixYuvLvVrgfrCuoAxyZa8G0lh3CSru0l80+8nLN
yNrj4tticLPFyb6/f6tuhDqFaImN2H0ePEXqgadtciiOJqIHNZYgJLHfV0bEv49l9WWLaSsSJxVO
NbBDyNrQJNJuAvL7gKOvGyHMthiyU6fGDLDy/HrMqZ660uIGO2PnR2hZWg3RXE6XGsm+isL84MFn
m+X5n+NWOf25CgsFj+JgbN0y5r7pop1RCxoRNvZbFoGjWI/GCt/W9IQMeYC88FC0meBQbEhx/4ee
tJdHX+/+ezH+KcuyNc+iihVrSwMmdYUvdu6MI/lnNnPecSqx2JqOZIVcilSCY3uMQRYe/G2pFcGC
txsPhLAFkAAH+h5dA5C10yCMIfjR/KkjViIgYsp47dqmtzYJzcmXZfMta7a5iyVaSk7vD02urStl
B9Mb6WYPRkw/OAG+0iJGQGJdo+5dREw5tO2XZGHfHatBfdFbRMcSRz/vwLxWaUz9MvhSUFyfmKEr
RcGAt+i3mwY/GBtnILsxZyZgUcEwwLv6swiqGw4fludPeE015deYOC8wa2+C3o/3ZJTNloqLXTl4
fBHZppD+7GhRrfnIxeoJNGulCd6EU0ZaBBrr6QBX97mdcfSdlY0Ofu1RdDcy/BetOGgh4B615Vbi
0lwW6Uc3jFd/DV9CKL03JAfZWav6avwzt89njrz+KraAIVm2/xWZhW4gzS/PvykTX7RIojtPswAV
ZpH8cW7fQYXcTuPzpB+QSkcePuCQsfGpIhFFupuOlxSJc3eXXUP9+bXf5e00I8EzPzUSVJm+6aNL
DHElr5fbUxIFMMYHxC55+tns+2CFfNBR4lbNYEx0R6J/iAuIcBjeubgyiFrxhM2a89kGb9z7Sf36
dR+e48kt8oaJh8+4QGGpHf7IKiCiKH2UIMPx++z8ujDcVzWgLs4qmqvVjtrH2jnzUrhfJ2aW1wPA
G1iGaL8q/xBVhzOAQWjRa9lgd0YddqE6qVimFZ81Db2PJUO4RMvM7x9pmT4mkwyYkQ8obNlUdCd3
kZOh04TMv/RuWCT/5jWgGS3HeugoAXuIqDiC/m+hf7F9yqfzgh/vFEFzUYqaBWkjWk7FWWr4xM+A
Lv0/sA5Bhjhy5SLgW0W2TUBVxFx2TOMScGsM0Oi4zm9SPJQ+c8/NzXTFeS6Fz5SucpmSY7WH1FNl
UvMoboE0ucEsSd+x2MQS/un2LOLiWwPO4F9wu6vQ/Mxv6/Z+lloqkDnlP9lkopWseoW0/e66g8iq
/rEXk9tQ0UtdEVtKwUT/7NO7qYHJOSHoZwmSEI7j+DIAORtCcZMSADxsqKWicQFnd4JOb+G/YNdk
LMaqhffpNtDUtaeCDj67smwOz1TPLip15MS78CGpRkKvY3qC1LncxIv/j93DFwttj0pyNGM1KJDW
pXcfVXV6WLjDm8UCBz3BVoBjE5VGnL4BviLyy6IRr+0qIJI/tFIHiK8SuAwNu2jt+81gV8Fd0HNp
W8THjz8aeOG93C/i88NpKIHyc8VVfOxMN1/1e0JoUulg+G8RxVN3z8XMH1exy89qymJg2DJu+snf
8ICDzr9PsgF3LyVMBConppAQ7WS2rWr8J97TKLHDtA1kdlUIEXo6j7LtXJkBEIv9draGgznoB3dZ
BfR8WbZVEVyI9YkD/gOiS1angIbFW6JvQU6n+EIdpybvA6upAXTvnWOM9DxTtZuRg7PdNW92qkb/
X+WMOJfbM97Guh5qoO1dm+2YKaloXNfWLFHFYtWEGFL7Kv7Y0dBOECkca7m+6VZF41gCWusVEw/+
FPf0UmELRCFEj+NeLJFSFjN+6SwEHZArPVg3e/uRL8kA1FRGKNVKISM2FP3xelYyR7ZudQd8UeTw
SBaX92JU3okIaGMGVQ5pg+V6rrVf+tmb39jajvz1m0Q2+wy1dKDlT2eaGekPsFAFO+C08kLLs7SA
7u+oaFhmcCV7L82fixqbZvwLqxze3udKonGKHctbMZAkRpNhyBO0en3TUOaqakVMr34wrXZMf2y1
8tQ+ba/ZmkchxqWrdBvUa2sMZBFDjB1fcniWv8MaUeFJdkkqxecEMNY4VATOW6Kb6I1PzdREHFxd
mNwyj34KwgD1SURfnZQASGZcLluHseldiSfaJNUDhepCDmCmZTRjMq/EiuUFqVih0Wi9+pfyjLWR
kH4g0mxIx6Mvkx+RQ04MdJ9ZYUq8q4/zSkTpe7oroMJsZIl65t9TKkltRG/bNHz70h8+RQxNCFkg
0sC3tHED94E6X/Gtg2zBYioNufZnkKdT3N4nz8lz1GDkVtd2vjlQbfMuOLKafkuIeDR1tur+vzGK
CfV2gtApILEeGpkA4puwSC2WmqKoLrsmvpbOD+NrRoeekbslrbt6Ph4QCla6NqEaqKskHqvR6O6V
MSZSRZxBz0DZxnnwbVR+OkryAMUoT4tHYPPrpu3q5zUY04ft8VuJ0bK7wPZEUmxtEYK+FWDnSHXX
sj4UQzPQz/1uw6ZCnLrxhRQEEYCc13r/fimMAUbWsQKdGWoHr0uzeYLQU4UmeZnvFtcqd8NsQhbZ
IrOnAvQ2ah9qYWIfs9e2UqdH4YqGQf+8ovcXRYZaMbVu+nW74IRlTVVa6QFQKjpnmaiRxGzPm2j4
hsBMBWsFeFYm/XGbbzcotK4b9D8VyfWPO7hDo+GA9wpA9E2e0aqnisF8BpFm56Q4Zm4/JAO1/jYp
Jr7oPRaCg3maK1Jf1VJeCdTtT0Y67/GYgrc6WulaUNLNHLZwnUZbyW8n5uiCJ3wLom8bSMd5knF6
wXgga7i8dZ+jomef5hS7jx4/n7EoEr0VgohfNFmRQjSihM0Z/L/+azbyhORau2trPI8g/eOJk5xp
JhrKR195hln3w2lYeGf5g/oDi/AcxUafmvNni5gAjvj/f+HPAl9TtOv8D56hGtgM0MkGbZ6nuoDp
9eoxmwoz9F4pX/1HPGmvjTos6jUP4a+xGmBUDyWM1Lt1oyj14y3NhNQPZIlluz/KD9UdfC3xDqIC
FqFLPknCsmJHUUqZtEwsA9wXZCRxhV+s7ZyUzztu7f00phWjrA9sSkK+UmyJnQb590Dl5Z7czBk7
M83MaukHBgutMBlZq0wJPp+V3bOPqPy7AE/KOtJynmOItyYvgzGLwe7PuC132wZJCIo0ALvQxd0U
D+JHmDEZsc8DSF5Nrk74V9MggbyvFlK0H3hF4CpvB5YIEqc8QTRjJf5901OXJR4MICn3KuJS1bN+
DmbLI/i266ErwWqxf0F/7FshHtnvJSWhb2AiEVRV57BRIMVnK1Les0QtRbGeoobylcMfi7QWP485
eKJydiXNVPt85Bv7cn2hNa04rT7y0bUyJj3n/b6ifvKcPQCHf8cYznpy3s/cauIr/IvnRuJi9RK6
qpeTCZz2SsI4lqtwKKLR490g2aBiui9J3Tl/GjSN96gePKUt4CVq+mltHS26ENIo0+cNCiEe0c6Q
WZVJuYqVGibb8F9HXK1TT+V9OEWlMjvCtkcFjIu5i5YiVzICYD63RRRuoLWKfw3bf0PEktNrXmP8
B9USDBo+7ct0imLcuWKruxdJNSA+ib3OvshmXZSsRlf2JGlSJ5llDrVg2BHw+9SRfKgV161MOukb
ISxwHVPVDxOGEiwhLkdZtVl56Ncg3mDIIrofF3BZpG+q3IlL2vJc35UTIrl3z+6hyN9AU8GLZijW
hOMc7h5qCEfkqg6pFfWF8fE19jH7Ew1CoXfeXztH2gR5KPVaOguE8XtKgZfvlQ5p03JuOuLVtooO
V/Q2BDkO+q3XxbkBq3DCEV7XDoWwjIwzAfxa6cWqMgrNpMIKTFjC8RxFj21JxmxLa0d3T8U/wG7n
ztDsc9oxszm57henVAWgG3Ib8YQklXt2PMrX2Tmsrdm6hkNUuCKTGFUgR9RMBJt5rsThDW48Yd9F
3g4l4iqrh5KYoYk9JMyxVa1sL4xJcG2+51o1tbzDisatZvbcHTiwdE1gelXL5eh2zw0MeBOwPlKy
kDyauSqpqrkLsvIYM0lPhy78b3RBWBX3pQggTXk2Svp4vhAdnfsaj2KHqCKZbw+IJqmAedHZ/1vr
h8PiE9U0sMbrlTLtvN2K9SDSB4I1uVNp/KhwurklfZRmbYI/aJhE3WjFMkBDk/P01xoW/YCeN1AR
gPQAEaa09QoRKzx67+zW3nZHsVd8SUdOkMhksjtjF5GhZL+TzUXgNzTijKzT7ZCnsONPVuKlIQwz
MuBE8+YxCf9T8qUUrhEeIrce1u2knB3yZ7dm/B16dMsfUtk0PKMyOQG5OPhPMXsU9idREDCWBXlt
JRp/8DBdbaF/dybU762mB9gKaUym72j0FYNUwJ776chSLiALOrgJ3N0Afz9SrsiOqdBZfpPojWfb
DQD6w5h/06JjlZB2Rl/M7mL3073cO2IOU61SMjoKHfWAnnvRAxKPakFNlfgQnmekvnpTB8B9BCTj
q2UPYFpmSNdW25urh0nlwZb9002fBblgIR6+rrBPLSCurERetvo2cMDKxfQagErZpBPefsYD6Rk2
tSQ5nYKVWitVG4RUrZlftQ4E/2nEugSphN6JEabf+Qheq5njA8c3UGF3gazms7N2GX5DUuAjgRG6
x9M/VWB/CMtEAZV+GxLeK/LfGRn0F89uS6Ti8HzXhuVqoaz9VnnoW3lmJQB5Q9MN8WI1skZT59Y6
XOj7qK3N4Z2IuYUTHRuhe5wQ3BP5m0XR7d9pz6KG3HJi64VdsVnWtEbdl3wR17fFoH/RD6rwd9/C
1JYwu9y4xVrEZlSwTivo/NG0WuWbwaAxJKb/TbauhIigKagRW0kQLHu2YqhMCMrQXBBlogcM/TPD
djUhNuSZV1xOFC2619FMAWarYXwelLWmUkZVfK8yYB71auWfMh9gKewGmhPaIDNHBZskR+q9wL89
Qxu0rrsgsgbeuLt0exGWX7VPcQiPizPwOKqj9NLTtrxejolu+86kjFlhxSbEDSgyuHcpC6Tc634m
PhBvhlgELj5fIGO4scNToZt/y+lJn9Zbnjvqws1bYbrP52pvwCK/8EySq55MfbKEF+9UJOOSSUGa
OE5Vpv5kFJN2XmIYCEY0m7auYMBAxDg2Wyu2mpS633f82O1C/haQyVmjz9PIf4ad8WxsIndpRE3T
UfG1VLAuLMfpzJAHBxvmOau3t87nydfPe0Xot1Dnc5vXqkKpu0Ymxc3TvqYpjXuFe83s22gHBV8E
kcSSpR9HaaYhTdYtdfz6UtumIBt7OxLA4NoSmdfTd1TcIUcVr1vsVVa1VM0CRoiXEv+aV4IOJuJK
QVEKSa21ouF4gMH1J0DWtvidInIdu5f05KO7//tVFVwi9zaSciW9AoFrKL4wKrhThvf1uNFpSn3M
/KcLUVlbAOyvMhdSKiIu8T8xhcqR7DBbDEYj5RxPcUMB4nPgKeFCFe3LbkhW1bqBYZxoY+BG5Df/
djuPWlbGohjObQvcZOXNOIDZWBEQHJsRDtvOPcdf2ikYdfg3DGW8Udhi+QY7lDQXZq9NoSetEeqG
jk2V7q0tQTqwW0xx97a9Kn3dKRDAToc4hl/QAQxAmRubZFDAZ5KiAkuvlu36JlWbEieT6WNZJ6gG
ms45HexcEz1HMGBWaLlUX3NgHqnzx/BEohScUbPvKSO/t/egwp87T1SKbz7nvvnFZJaVgkBiqamU
7NJ27aKI/M3pjjrbP/YKYdyvIi+itsKFG1qYm23TTVyYtERWl2g6b/ykv6QzJyFsG+KQ04XNc7sd
8W186loqesFD4a0WEtHqKRkFDjZhdj5ffcWU3XVqCgFMKPvfVowvs6AXqUDOsNtWZEmXYtTp5CTG
iHqpcMwvM5IoQfYH6niWkKQNIVYDUu19VEoXuimm3UFAv0j18sHKaHYi0Bqh52iaMUMN0NAqyk07
iByM0FUIp3Q1POjn3IYKxlLwrLxU9W9wcUdKCrIyGJEhfccfnwBrOUy/wK2OM7irir0yrvrOvlzL
hW5e8vEAa2buQ4C6f4uol+uspLjdGVz5axBvivPFJ4HEuF1kWtJS6FYh3u2bORbA78TUfnyNfSKI
pp1zEGQHYOA/GNHy847fgtO9nR9f3vvX+CKG5WE0JWQ9kA1RLFKcFrFYMQmTL7DJhtgKrlF76CWt
0hAhPL2EHk8n5W3wmPPDAmHC6FxLNmQiLHbsXSB/JqRbYoL1Ydk81aiRRx6lz0NOsgggtuBsUOeI
7y5o0ZbxhCMb16cup1khq9s87WVPuCU8pd1z74j0YZlo5YqQWshUTSoyqx3Kh9BO5zIBNazdl/Di
0PUOqfJtJmIWmyADa4hKY4Mlu1VRD+brLKulLImPvzJpV0VzYiChhjt3YMOLs/w6SGEYDDlbbBD5
CJ7hNpqQ7vQZMfC5Sa0iNFjs6LQfYN+KFWUwmW38kkFF5pUS3iC6iDAwjp2/SmJFth3ITA9Jo/Bz
4DvPxgPmqt4dpt4Odu5wiV+epx/ztyBcQvgaob7r2KlQZ68xlGR53RmzvRsTMc1/djKhThAEJd75
FrczE76MXoPj0aV54+ctsNAJwabXZyA7baBwKTJi/t+JmM9axqOkQ9RiFmEce7CjvUVpLmSPH54J
9/a43TF7x2hyuyQUMyNHA+EZ5/J/HLID/D8s78YUTu72iDJYxyBkCkxOSN62vbgDjuJ6ZnBopF3j
EoJkLClVNZ00CYHpxyIynciTzY4otgYb3Slb1ED3CV8coScSAqB8Rl7zQB5Er9q1IsMB8hx5+AJp
nSgom3Xo0IVt6wDPh6m+skhHuNzEbJft3jNvDugl6ntffOjLSS62XBgLE9fk3y4HFTq7splvaIK7
nBFrRcPN4bsDZXFKuYQE78eh/iUyhc1RieaQedn4I9VcOXNEzJ3q/lz6TWdPff9Xep4kAZ4v4CeU
J85fXDnEiXgmzrXrJ90Coe7DGZT5dt08lzPeFmnVxsM9WZIfzf1z8aTZQgy+KctCnLA83AjsE+P/
qS2h6EuUWLokYccqzyhznApf7rDpanh3hcZSPYHvNg1NuA1AZnAgOseXTxl8tvKHL4udcXR1K9oh
HH9Zf0mJsE5owqkFBgh0pDCmpx/EXb1LcJq3NXMwvIV4z3OdXu12Nm61Nn6hzVfyl/ILCCewmDwc
Ho+9Ut2n2prHMun18L7NKZmEHaWboTr8h/qKlP7T+OChMw9cP2m3U4VEvyW9PNJDFz5mATmnIt4z
MoYE/zZ7wgx5vkAAcrV9cElETSZw83T9HdhN+u/VEQuRTGjCR4d1tCgEnU1bwufV46FJ6p2fYO2Z
LPMKyU2QhO5nkEQ/R0KQ/WIobOuihKSiTIrW6mQn5aBgDgAH+JJFgBqN52YQVXE1I/S/FWKwDYvh
KTiKdDYG6JvFcO74tiWkEHXupRjAJp8fkWg3lUYg//TwJlfoZz03d0MG6XEcocHaJCO4+AJSX+24
xN8vkElmCwmtDQo61DiFi3vqNjM4jHfEqwmMRNacPqrRXMcqvMXcI8kk0N0oOU0vkzm7fQF/U7kA
2dOLM/CT8ldf49p+t0ti5pWvjGsn3CDtMM+9UqYypjJT/EQIspkqmyuphBaB4HDlrb18NFrJgei1
0WrI8Fs5KjvFX/cejBWlVW8XrXCkfKRTDsq3XHTk0JjmSHlqsBnmcFlv94iu+y36oGJZ9ZHmbpLI
BacI88MdjpWyphRVHOivh2Zuxy2cDZ4+upzFxhkL6rHcemTh2JqLK0LDc+eg2VNpzTTfT79pVVzd
YcRb5+BS2hrLiHFoylx3BsFgdqbsUrONaYTKEG1sqR7JDKmYqVs/xQP5NkSnu6i5tL7B8lBNB7Kl
a9GuPJBVQBsx07+94qFr7+mlQIsJl6a3TQeANOvQqbxQ8AbJknIczRkQRuFFwiC1DaqxLMo0dNqb
E4W5RlGn8kIA1CQy4rMYRIgOBoFckc2mq7/QznqXy8Y95kv+jo1Neql32nhYC5vMPUyqRQfRLV8w
XAfVxojpIKIDrXvm5VlioYAOj1qGJ9DsBV+yx49ZIczYHCVUO78nskgyJrrW+30uz+yH9RwhOFAM
PGLbG0O41jGwRdeg8i41kfL2NbyxqsUUFFu0gQIsUh2XnDhIjerOGCyYNN7sjKm5gzfAFNMDx9/z
vJK9ltBFPwO2p89ni4V+eotzyD19O5sqsO2KTaSXryGiOR/L48A/hfN6ADJrZ2+2k16jl/gGawiW
bGG7LDfw1im4sJtXdmcV0BNnZG8VhdS0ZL2WaMCTmOiGS5GmvXdPHuFAJ2GMa0jt9kz9UxEyAKM9
F2hK4c0bf3toKtKr+2ySq3s5kfKpe5udacjn3k8i9o3+D4ocMf8Se1gZu0KlFwqL5/zxiRr9MUti
T4c/sag44UGmNZ8CtU2pds9xTY8DCZA9VxnR0P9xZqlL4RcM9V2dVu+MgEPE9Z5dAY6V9FfWHxhG
GyiF4BU2JKj9CsNkjPE+MiR0WLivZXBmIhTv0boknTAWvpfdmfF8F52yZdl4x3/nLKNKVADJLK27
bBY59ODfbG6TQgT4VVra94DM+YEZj5LjfNj9/zyeHAdBirPCy8qfvhXtEQvDKI6PrzxgNwhOW6Gj
QLwuNnKWQ9Ouo1tREfUMctrpcByG761oz3cbchAen8REcsGBe5ncovkkX7CFjI1MWu3JZ4Ger+KP
f/u31RihnlALAHwNacHozRA0WsnDnk05x2iN20YtPvGN5JUQgSomDMWy7d2HQzP5Gllh61f+UIAp
1hi47eRVLj97CfWrwNw82kqcHfI2oi25ZKAe+tQfYbWLI5aWQ3DQSuaveP9dQBIcd6D1RpbJ1K/X
VJleMnCTcHPlZTlhb4wsAKutudNV0hnM1fnL9cCHyzKZnXsLTpzomw87Tgg00gqgYwf5vfeYGQwB
zilPLD3UKPgX0iWUHqmzHdnVgUyw4fIJzoMo2BZIEbwGMSgDDCnZ3jAHzat+Lh4LaTYsJYwd/adQ
d54kBg26bclV5gV0b7C9GBwJvH2qEjaevY7jMrWKORpXi4l1HJb38NctegX+QLOz7mjs3xW1b8KO
78xo3s1/G9cUD/WzVx/9FQSp9YS7E27gqD0wPQjuDOVztpHQFp+B0ZTnw08muO4yUtiluO6Cr++K
JxDqhwivJcMwW3OvxdAyRmGIIt3APK7OnG1hAipMRbKUv02Qi72aXLd659nE4UDJyBv9t35jQDJE
BZ7eC/vys2IzuMrrK/QToulRGRoDZXs9ceEPOsFFzduPFEpVEP2CAoMROrLgDbYWl6A3/jQ3k5pr
1JsCtjBYQMrR4dmwkN8oCXUX6ougHJvIGk6Zn0pu7HglG8T9D1QVP9gCeVv9UmDzy4HjwMiEGrw/
f4n2Qxc8nt4q10oyR2vt4ua4xv140g7QkI59T4Do/5BVFafXb82agaFLor74DT0dWKnZ9parGKBS
s4yikkMyyRxVw5m0nr5ofMrk/EyT7d9HxOa77DQm62PLmnZu5MIs6vRGf+NjaS2BDlhCUcf2wbOa
WAaPqck9IyZYFY3IJQelhwu2K9VJk4YiOrFLY+6xK0z+gCUh9FfCb91VhmihITp/RYL9a+g1fMsL
kYuQoJHmfE58Hw4/Zt9aguxWYWTId8tNVTjXZs3KuH39EI8lPDO8qqBk501XHG/M9zH+fs3VO/DQ
GiaQfdlpV30isjT3uQVQV2vNIQp5xh3xrlWJTktlkXdc58Sg//nOi6pLDnsmz6ZNM3UigUxKXxRH
stsQ1gGzC3OQZeVcbdw/dqd+I868inhCpe0rplIv5vQjBgeS7JqQjyHI1cdxpu94C06rRU/Zg2Y0
a20hp9oX21WHhgYeo8h4f3RTrJw5LpyUwy0t6VUqsmcK1O4zxtsZ05+14UXL/ACZaENpNo1cfkCf
/maMPE4qSDt8Mg1BqR+lcuF1fXg08l7zxDysY0oZzMXssZ/gsua2U9V93DR/uTsPt3Fn44u2dmxh
r3zmtc2TA4trOU7HcFF6ARGQFE9r/2xQaqH/HQJWmDsn4xyQL0SZb45rVezUl9UhPO4O9r5UcqlT
Ba67ZGpGDLgK7mkggdSRRF47vFe+2M89BYJ/uZs4f740FywgDzTJmZg7IkYaAs3s22WFtkf5GsaS
K3yogd2oCc1jaWhkK5k1jwOcT7xmqYIx3kzEYosOfdJSD0wueqZwSFK4LjvXrXjGNYQtbn5yK+R4
YjSXuX3qWj4YA/CfDgZ/Ytcr/HP7cGAyzmloswpQmm3/vdWPUrlPszzA+s0b6Yv8GPioZTTYGBIN
boEdzgsBwhn+KPcWqU67noW9VTMjJ3sTj2f/Ik93XM8KEQd5Q7ymJwHgARMIfQ5C+mGczAJAp+x0
2gtTC9MmgkQdWAq4v2De7HeZPQs0dqJjtSQ9ID3QsjmVo6locMGN1ZxoMCg91wCwQtrdtciOyAuk
ijJv3o1nO61oUM72hgmh3QObNPc4nDtYDRZ2Rz9QJudtUzYizpiTs7i0xqFxfX6LKSzGhG9rFvtU
/TUgRWjbRnR1T7JZq1/nq3HE/bDBA3PWpxmbs2qU8BXa0q1Sky9whdfqKfCqK51vpP1u0jJ8IdK+
TICUSyN7mmxSoIV5lgtCX6q4ThTo4df9hliNC1clxKXIAd1DAdONn5zKJBNKJJXW7O+N4fKb3N5J
M8ln5DLcpZMC2q6UdValaenyZFHzHf317ESZeBtOG+2fkbuI8aolXe5djQkGt1cHCG1PbkYhvUhi
CXx3DxJQk+R20ZLiK4bsWzmxaZSF4Oi9doE4cmEpioy+8cVnmkLmlTqfMCYq3g5q5bLpV+lSqEal
VAMkcXf1LGFuj1FmlCMiEGogl/sKqq9YIkwIFQpJV7a4WDHJs2ePFD/VkxvMQSCh7Pn2/ej9GyjU
GHP+fnx8Iazm8itwPKpUT3gLt18nXFLVxAC9eR9DVSliqn5wX+xoMQn2t47VVsTl33+r65Ld4V/J
mhi9cOOMKIKu86Omy08HUI5TgE2B+dxyH4+QyH0Ymx48ZnDD1DL8Pvz6IV8C0f6l5jy9Mi4zSYxW
p0siwUsGTmCNOeq/DfeUjeMixmVrEJXcraGSvSqKe8DgXl1skZhH3I2pQhuNlYJGoA1Xh/Rwf7g1
1mQb8ZR2pMKg8NbKcohqtCt5edxBqmpTTz04G0yR17TLGIhfPOZQ9T0RLm2BnsnDSTQPASLRlNph
rRVxdi4c17eyYmEMywc/s68DsTkNSSs5udkJwpmoQfjxDc+AAFoNEyfcfz9vrGCmgg38FFyFmxA6
S8aZpBv1pwDGRYcGjgA+xyeM2OpikZVfkuj2WyPVMBZdV/dUt2EKyi5TtZpk2CMW40Zw/0xqMErk
FuPkVTcU37abEd9yj0/sfjhOJcY0IbzYAwG/sbJIvxR+jkhAjFUIX35TQtmWCNevDmUg6YfN3JvH
M/kdIxhSwjJeEbRNssKX8nunyl6rR2+/bkIg7GuUri88mIhaW1ftdglcgAqgmWwRT7yjIls+9YP8
Wl0JSeBaDbSQonm8bFZ+C9X95lb9BdAuhx7uny8lE8onOiK0g7Xc8BsgiOiZT76DG6Y7bXFUnqSH
T44/deWzuXl5WV1gvxs4umTxMTjzps7+uh2nCmQLCKwMrC9WBDjXtzs20ThFx4UWacjI9ZYrfxfA
bI+P2ZejIwz2etQbi+H6SsZlG/O0DEyJw+yQqd4u0G0xKST4lIRr0UBAnLcpJoridvlAF+zoRhj5
nTEpYqlhm67YTXrcbiQ88gJQ2GXo3amR1l5/zPoRX22JD4dLLK3krONejdwlKChw9xEkAZI0M6Sd
LdW0bKgBw7LhSY5rj1DQz9QZx55dlMdYzvJaDfQpkRMkDX7howavVFCXhZwKltu5Ke7MrOd5wMRm
5odWeLLCFKWXDm9RxlWgsb5vZ1m9J6xi/hAkrzgtBRfcBy4lKD/JfCMfg7XmSz4O06eg5cOsUBP2
YvApqflNOgzcWyW85xTKPtOBp6/otZQP2RkiGXUFc2widMYprL91gKs/1mdlvmkyd+hTaNdaf2Kd
18d3JfePhgUHUlfANzfn2+lKjCSoV72cHBmI4J4tJnbvV8Z2JwG6PqV20l5FzKfsvJzG2W34+/tz
AgGFQMpiM3oNZpzMU82ZEtWS0WZ1XZuSBYYcNl5Fue9HkC40oesuVU0Teu9d6cQIYEs8tntDuVxa
1LHFbH3TvPXV2GClgfdvOlGVbfJwDktlc3dN6em/vOtBVwIkAgP7I1n6TNisxWOvJFydIg7qBQl2
A50zuz1b/S7DAiM9+ZFm0IOPg6J0wvaK8nnMmJ31l9rvwCWwAvkBc4xIlOVnOsyorJ9lajnD+mie
dVa7npCyoPhbEDwgS+mEIAQGH1uC+wLYb2VDDpRXGAxurmZIbobKzQmEB7OMntKUQVy0Ozg9xDMq
DyvHIRmac7XNDJQmbiIlvZBsfJQWQ0A4wVh7fnAlMXlO9v1azl+oB587T7EPphOh4MS/vPYX1EAK
t0R3K01WOinXGBzvnA2AhmZ56pZ9Ftd8PIyIPJ8ISuXV1ENMnpULKqzTt0TFML/jEnb2TJLBZnxP
NCb7lIErzECORcQI1aTXYa3Ln1NpUg0Rg/Yslu8jFFH3HU1W1h+LG8Ed3n8/+jkbFSavvhaKZW9B
O1gqnNztG48c7ALpK44sgTD9amVMsRLxKTLCbSHXC+qBTiu5OO75Au8+IzROnSDDa1rN8dwU4+no
Uk5DiCLnF6FQTjJUR5lK/aY35kWxf3lXDgHpyKXn8OWr2rwWr13D3TVKco2vStQKkRyCxNTTuDzb
yzI5+SD2PvZzzfnQIeaz12xStkHjSV4wEZwjreynpFZqYX+z4po7zjn46hzuvV6hg/gORBWGKila
3ckpbllDGG2FgOaEmxzuXFgHd/W6tln0b/ySoygh5k5gamfG77kwZ1K6w9sK1Bo9I9muBr1wfxzQ
qrQ84Ev1/G3gBdsEQTZ7kfr67QU4ICv8Hyl83/w9Hj0TgAOPndprSlJi2tIxQ14PJhdTnwlr9d9S
U4c3yAbCH8IMqtFiMN3Js+FTcavKGg2E/07cKx9QjKDOwALm3UZOSVwVSTVGC6Qtr4J0LbVsRwyw
BabEGvbaY/pUCdrjkY2Ad0HR4G0LApJUW0KOm5I/vseYGyOo3W3Fy77mdgZNKZkKbs96xkdOqtzw
essLMGqz+4CSFOaO5ptmhZQyIZJ0b2W1bQDie0Q9kUmZ7NhDUKaayTmBati3cOZFb+qu/HQOhjZL
+KI8xXnlAlSe+ugoJ+Lb4FRyhUPGbldcPtwDbDzYhJqlCi4Lfp1EHq/LHKNvynbRfSVFHa8F1+Ix
9f5qFJLvhos+PeXoFB7h8MUK1hDXgr23gBuTr7XPpID2CbjOpo76G5GaLVS6DWvnAA92puEQ1SxH
DMRK1bhz6CBUUPurqRVBCeN1onXug6M37Xp9CKfowiKNJUFOnfIrWfCvNqwdpivkzmXlT7mnEkRZ
JiER5IVsunjs3rTQWDQyq/qAyNk4Vk80PujqcmplI1HVesofrOD/4tNibHBQRy0dayH6Q/IpzZHK
wgqnJBql01+M7lsyW1IOu4Gs2GxIQv9mhqkEdoIHdpwGoUxMjwKRbWthNubBoqLUu80RvfQCxmxJ
nhKDN7kawJcoynfHjfk2nWOgQJZ9XCiJAy8uRen1pcSXQ84nWWgqz2MobtF2PljlCA5eYZugJyRo
/2Nu5J9tTWCLXA9DgVXtDechwMkDRwQrYJd/vnthhlfoVZf/XpslIcQwolpznhw0OZCbtiZqZMFT
G3YCVf99jSlaXEB2i7oIVFFBrgDBF+AMVIMOOQJ5dVNy1NEht0AdfqTtEyQ8zYqQotR5Jv3fENRr
zWD0X/9z9gJlLclWl/SQ5FKewDerY63pedoLb4djbkjShJ9uIk6gdjcPp/OsAXrbW/KCxA6AIJb/
bGR6CcsaRbgCLkjcqQLZt47S3/3MBhhUgmZ37cDa3ICqVkSNkTy78bV/fiUplSREUi/3uYPeZFYQ
jfIyRgIeHLjls4TsXu/+aH5ObAmpi/+gk9GHftPjW6o7B7zKVnH8rR7tn1ZDXLsqm66vjf8/ZO1R
y2fapS7XWOzahrGbVPZIzeLJAwpaVdTHdv9uu8OH0Ol0Y7mtU1ka/FyBFOTSm7cVJiawyLwz31k1
HO7IZSkB29kZqRN61iCScuRFMRyKzbKihCscyvCFlborQyLjuaSEtZfobvtjGJzr2Yu3irwOneT4
g7aYvlPzOMUJzNUH4sxaExQjVuwT/CV6fWN5vT626IWL6vSci0BSdEpMT8AOjA0AtDSIgFkp0HX/
scwW/xV378nNg32St9NKaH8SCq6SFT1pLitEhmj3a2wdKpG0p5jLLn5tAannEBZceqevPyuLMSnq
b6DBugCu1D3SAwaSMQv4N3Qb0Zbx9gsUjy/Am+10fo3Nyvz0witbJASJS8MPB8tb2xgEOFZNpNWw
BPHa1c6CctgyJt+V6+Anb3ceY/Gfz9sd3sJCOpMZvdlxk7Qyto8ytYgsXj13mRrwxV18qM+77ZrN
iwdaiTizfY9sn5HRYoyFsFAoXpCiZglns0txHL9I+V6k6MPa/8qoU4HjKvyhVeZFU/Ab5M2EE7ry
3veVeQy8/g+E539eCQHJ+x0E1Kckjde4HiYCVuFVmGOM0ZQm1xkKjgA41kd+MbUGej1pN5FeKGiY
7VffTm0L7d4EwFYjetaKawFS9fNo+FbI5XkYEfhJdxOqcU+meRHiqRvSjsu9AcixHpBQ0VKYl6cg
8I7pVV4FjmCJ10MOREddCP4ZCgvDChFKU0eopS7X4B9f3Ji3+sPSEMsj43V0c8k/EK0DDkZdxTJk
LLQkMoAUFDth4LgBVXp1I9x6B2pvXQNVYXEHYgkcjN52phfl3n/vJCkagHeiZT0qqiUMus7m36s4
ERqwX831R2nonyBka21OyjjKaupy4BVEIFVp4BcJYE09D5nU+lBmWbU3Do2bJeXqJfG/CkUI9qLe
iMm++SHofahyvPjzN0oCtaLncYJs56/6qoge+Qm7KezYyqlNNvrj9ku8vYwaC7sLTPc0jw4oNbLI
0gWAbbi/nMZcc2q+UbO+XS4QqUl7TSJK6HqGn10nnwF+fNgzLZA+gQNSXbdu1j2OTft8WnY6JOVL
hyg/5/CgAQHFylsRwN0H5ZebAsVUjWqdKILuVW/G5uyozQlSDdIU5YHQEYGRuKVqTO2MgEOeWYPI
1gBdZ4TylsNqNJNWN2Kf2ICyUtWY8c/ki/nLwbcTkSmIVxHMOj9S7YSLXmDQW5oqjaJxwe38SjBU
oZ6/1cmtoYEQF6sxUg3GvT1bj4Msvw5LeApcffoA3dlZ6HUtgYCv8Wj9JOklOB87Xue8N+HyljOB
5/R45JkJM3soyIsNCxLTwmSUfDNKVCID0S6yn+UJeVQuST2YYm1oVLR/MRILZ27Xbkw6x+SBKV7J
fP4JpgC7Qc7b8d9nK/T+3DpW7YRgQyMgRlJ431gOb+onmXyvZp+wjp5qKhDbPhQshDzZdA9DF0sc
v0ZQBzH65D3uCT3nPWJ/uFvSULQ7zs123WUm+NyPcLw5Syh7NX8HVrvZa6MGyaFNkWpJrKr0e3zp
lbvN/AxgjJ1ZGXUu0PNxfIieDOHoeT1r7HofKl+Xll+0J4mgfMFeirL2sWfw+A+BRK2quNHzNRyo
Nj8/NYXIeI9uPhf+qT6iZOFm2r2l5Z4qOAg0MNWaF8st9g92LZbLIUcka32RinGwT3E2yVT3mm4O
WMbCejIgCA+9YeXwC8/tKu8Qwd2kg/+4pc5LGVGBUiOvOcmIPZuFV8Jp9OZD/LpVyjqSwihr0Vwx
Jj+3yNPDNwKm2tgK2Y1xARDLYPpwTYBCnmCnXiyKcas2hEFWGHNic09Of0juvHoj6QJz9aQttghk
MPeI/54PMFBmZSuKXJkml2Ogg7X/tbE965lLYTaJBe6zubyD/P3URnUgNC6B3G3I1WdOJH7vCChF
Ry8J2anC0xFk5alJV8+ivLX3vuzrI620JjAxYSVFBFWqL297pCGOLml6bR+BEe4tzHDNhPL7cUra
sAkd2OFuPFKw8FHSMsJD83OtgwZja5sQnQPOACIHL+f2wvrsMqazS5e6ulfHwsIgDgITYcF5BL1U
0HSceGi4SxI040s9cvAP5BZHue4NUti3lotpSbK+PeX/qalWrbJlPartnKgV0rndGEjVtr/XZf/f
3+OuFF12on4YcR3sW9JRYaPFyK7hywslmoLHuAc5ft9wwdMxuNex4WPKQnR5x6zSGU/o3/Kkla07
p0axSOkqMBdVMu2GolmTXvDjcOqFt/kLBQ3u99TZl2eN/ZHPj5982eEQ9FoR6+XyAWKoUKTRVrvu
BreRrWMIDCiaJ07vMv8R00ctVE0bIuTAMgI9FuZ4JLfxZGemJO4TkMdmSyRE2lsu+jNPsPXzf5g7
mPcFpLp/b5z6reDWt5q8lqICCBie4ym9Ithwebp78tBM15T5NCEecro5KbhDHQNGZQZIp419OF4P
ftsM14i+F5GntwIjedLnTzugXspM5ob3Ov0S93g/lPMre9jf6AGnWcKja3ct0fAXyls07yjcPm8c
FdcRcQqmwzxAaGBCS6fJP/u8lJXjfSEpg4vcnUkKVBin8Omp8m+42/r3wWiyTOZxR/gOM5HrL132
Y0z+efshh91chEtGSusi/MYXgS+5zuNyWR8lcQRwaSS9lhsAOV8txy0/UPOP7NjE012wA+0K62Ci
hCSXczAT//cS85nF7Z3Miphw/7onbOEmJsnKoq1VonibQ3/1+ttB5wGqbqITxNi49bU8Gl5vxT/a
T1GEVuh7RKGyHH8dOqhqYkyPR7vaiFljncad46sWHPyHvrfXrOD1SBh0Lpzcbzw9/erTvVp5sPyp
KkrcJB7QPsKBAgO1mPsrTFzssPM7LwPa3ymUgulwIMaDO6r1ipv4yUlvz3WaCxtQaO/vWxUmd6yn
uOVJBttqHHwABYUNLgZXTz3UIGOs5ZAo6nI2PH1teDAPaBOmN/E8pWUfRapVw9qW24tdNHtYCmlc
guDplXMwzq3Vm1gv+RM3laQAQceag5xKsYOShietvM6/eBqH9rBHjT1aUmTWXVReQeoIZzB0/CpG
AufLory7rr+6F3Rc52OwU/T+TfA5i0qHqsb65i82UU21fb6H6sn9yxvx1huEJgvwH37unMjpiCNa
AGb5Yi0in4ykla5giojb0qwhWTzBoIskN2KegxYYHAKL/n9hWX01rO5lRMTrXURzGwT6f0C0B8/4
bnJUh1AnTWdO05kPbHm56jZZqA7srF2YxxAaaTz1Q+lJjrTC3ADX+Swg6bej2J+i/P9+5p7qe/T6
XgFLlnbV4NyUjHl77c8SSbFe7LyRKuCtqZnqwWEZCnKuFAbF5E2yg5RLUP2q021h+5Bf0nt1NVlD
VmulOA/stpQENq8K9Su1LO5U5kyvdRhZ6HDkGJZUyuC1pGiUPjHVudspTgg2SDV5ktbWaVKgwclL
M0GSwoVt2MIVId8ybc9Ib3O+Fql3wOyFWhep2iOC3fKlwsIXoBoVcT/eJWJtFvgG/5yUIAG8pt9I
Qg8ayCc3Y2tb9PO8dzMv+o+TwhS6cevYUz6YbnCTq9XWkt2TJ6UC/ZDgN5g6E08C0GBLUtSpfKqN
xxTwstPse9aHS/7lc209m9l6ZOdILN7A0Z+PUcTVNe+2HJb2awvc6PAYYnIOsFmcGtMsLjHBob5p
VI4PfOhbL8aTAGKpT+GCi2iD+IeeiOB2Fpt0+xX78yA9l1vqvNXt6ufmtK7L3XpscFlI2j6f/D7Q
mLO9sbJrfr4sNjnGSjwi6clwuG8Ae+5p6qhxky0g+BLCv6xt3OYw28RSNWL69GvN/kC2cCiYmNOp
sttVMtvrMjR19yYFm0XxkPi7VfP2LeDt3sDdgvJkeaKCuANBiLO7114/R8ukdJPr6VPYADUEgSdH
nG5P9Yq9/MHr8iW2QR5xyjVwVlrTfSvcjD+yTFfkg33MdvxF2RYBn/LsHFT4gXTQ2ZD+DP54vzx0
UOF/lfe8/Wk7GYJ9DpJrMUgNM1Yhc6HxkLDxTEroXgnRriTpLOyvuzpWnMt13ZXVvZKRsSSpOph3
qdf1t6h3NtFyaTK5jeYynNy8lHmN0GyXsnI+albub5bRhowl6QqCG77eM+o/gr6mWMBDHl712K4d
N2XU/mWU3VIHcFwU1ccR3x6/TmLH256SlsVHoE9EmVZ3CpSV5tDv5w9M74Zu3pE9slXK1AiYtfV9
rHBTIjKkmBhPRbOXKAaRsGyjzRcKo1KzoLFMW+mo4q1umOWem8vcFJhuWbeD9P+ui0wCN35WJjPy
eIqV8Bda+B5/kWqkxfJdcuWiILfXWRPBbWtQ+Jc7KuTAlZBlwCyTzT2R5kIsvxMPDpmpgx4K3ubs
potymBpFVO6/kbwqpc3zXZxDXJ1c39ywuRGZMdpOxd2sBWhktEuAhrKSYNvV7ZyJyM9ks0k+Q8bT
hQnidnNVjoaYyZ6YhGyhdrrdgvc9L3/eLQxiMAxDxuPRgweGCinL/s+Vvgr4CBQGJvxvWizR87aw
o16w6HvWtZpzLo/pgqU5OTkiRJ7g/3sKXAk30ZnDmQ4H4QFCBuogwkwAeuQIVnPEQrG7EbIERVHA
JvpLvsziTUF5uxaARRq1z1MrzHKj5ETuIW8C3DF6729AZwImrei44NjKw+YKzN8RBraj3hGX8H42
V75aEdlNfvFkdEHRlpcD5aw7Wb6NSSEn49eJdye8awhSOkhIpjaK19OC+VSMG8Y4YDERFWq9p3Vn
FtEYCn+9O8BQN5k1ikiWlo89ZoXbnYjsvz/1/PIK5NzQpsSxGxEJkrxVLbDBE8MOOR437XEpr63a
ikNqEhpY70FjZRb/LVi+QFVKoOCOO+qPAtEFS7lV9jP5PTI0GjXoArlMEMSshI3euhZysYjF3XhC
+hlRD7EG7iQl9/bDNaAtT00j1M1FxK5Pbr+7Cq+yiMFhUVE8OSU+70hRJ5RWFGurCVpObE1WhwCg
THn1t45KcEQc+6Z5hDWig9+PYggixN853OjPiHEdcdPvJNe/b5C3jp3dQ8/U21WBDjwXWDAlOJWw
HJnayAiY8rXugULrT4t436mpM71dz8CarOrffVqz8aR/PqD+XYKmETW1iCwum5w/2OTJpKSaJgsK
/avP6HVuYBIW5B2u1+yLkoDe2o1fkSPOIIO9k2R1Iwu0l0CH892KPxm5hlrtpBfuwTpMObQ+dE/a
QsgmZGXSbYv48oBqe1xPKyWieGfr91jfwEJ2ESVFTPlSQp3QjQFz93AE/hhGLecTq61ufyLnTkJA
GzeKoGbXOynL/iTgh5dLPDIo3+lDa5QkMrlfhkexKApHRn7IERtN2oE0otgS12sz7NpAVHpsqr0i
g5PcL5PaoMT22+Oc7izKNOt+EtFXG8eEURKh+duIUEjFFHaAal5F/8xfBrm6UCKl+SADecQvGgRr
az7bBPDkoVX4eAbUrvMnZuk/v8TrfsfM59/dh74I+TUgQk2nkf7aCaQS/KDP78QiyRAsD1Vi/BSe
TT8EWCmJ1D5HOI/DeY2JGJ3pw9rvuMguEn8hA9wq55N2a2GTh0hawFFHjDf7IFwAeOgW22FSeXSJ
bc08nG2rVFtfysoFbjo5MRZs2pazZaAA2GGBFzTMXTeVyBRWjL+/ENyQflNCPNrh5lRLz2kvIyhE
3xFhzHQuPzLzWk5/IjTmGo1Fyg6h1ZdT6dz1B3fbKxD4ksLHFl6m2VgXCnkccy55aMLgeA7ZVk6G
0jsIPyjpiH3bq9+dYFIaGZbZ9TbBOxUVMCt3GLG+rvpZ7kjCYUqzRagpcsJRhlyYclq38xlW7bWd
WM6l4aC6CF4rjrtBHDDzmTOcjcomrN8IzvbwBrWloU+7UsMLkynmHv5iK4jgX0ZtYKOFj+S1dYuC
dDuYV8+yCqtrRWNaUSN3LDloCYUjB7kuHggZt56gdDNp2WDJalKXCcFgCs+vU/jqfFId4pBgSIuv
wwSSUJ2ao0QQGE7rVEdvGpG7O7rNlOnw6jIaBzUSc4g2L5FvIW/3O7Cps1gGRXu8A4kZ6Y5G5ARv
g3TVukTfJNpNvlb/wyqwrFI9HGeVle5Lu11PD8oZWVurExeBIfIcmfnpYukL423YJSaxMKGX0Nm/
3EErWPhl5MBGx86TDVB3hWMqcl2cV+ulO+gkChFD1ws3QgrgxWY3oSiD1xqX3e0Mf6pYEYTWTEXv
Zca4ByDPHj0BFlCF12Qi/mGN9IafPlrqjHR10JT14BcW26UKMXwZ+cpId/EmDrGnLWpQwX6PBu65
MV6tSBcD1j0DqoQp5E/q3iqdZdyuGm0CkQvKIXszPyna3eZdKfsqcjEREZsQfd51EV6a7LP9x4QG
TfQDVu8sPccbRjdYc9TaCc0ybqgDnQuJjDcF0UA4XOuILSo3SSzzPvoEZC74TfGLsy3BEXIjhObj
/JPufRx1/8f4spgFWo6GBOSCk6uQJNxA76Qnx8lmh7kpmGn8Z54nN5arXdSzghFYkshQvgg8fz+w
TZpBYwNTWplQjA7AiVaRCOh6yabx2aDRC66HJWtAwrb8SqDA6CUfIWfNHoi5NqAJY2t7ZKZRtOrG
Q7IUXe4msKW9uAsxNNd1Gful4uKfoTzJAtdtWq8axaThciXHoyrumMEkv3vmpKkxIoYxhDR9n54F
ic3YfADjww24gse6yKwiL47jamZ8H2SrtHh90s5dbiZruRwMWoAx8yUKbJQ+uvoBb6wqXoUcoXas
HhnC7WajjpBzi3YcEUIktprumZanS/fm4ffdgepmRcMcznjFj/IZKiPtq8d+Zv9jOviUyqZ6t+mZ
2rG1KXjyxeqzltGL/2HTKeZ5EnCQbK+i7zk/9Y6IMtnmc3Lg7/YU8Yx+HF5f9a1r4uR2Gy4fiqWv
7JZpH3rpz+RrkTLDbTWZrwgy6WWeigzu+UpJVdgN3sgy4TrSZkFC1TdzwzD0sW5KStGfqKGKVU8T
KUTfXxWpWJ3L5yHtdfEA/y1gowo7CbkLFH0FNMtouKa0KO57SsMLADzSoIiI/hsWOzoEypoySEkw
D0xL/fgLAfjJPlFeeVhUQKhWpRuBx54eNqKdCzx9cEp67xin8H7iUlFNdNrHJPoSFwX6HJoHywUZ
jb7+7DLVryLTRxqIe79g/njiIeRKtnbUSe6EvSYL2kuA1w/XzIojVnWvwSgnkWgA8ma+p/TmcDXk
t630vwiTtnSK25NbsVoxNO8z7DmuJRjwQ1B1SrEplsCZo5rCNc+RKZdN8aPJ+InmWiLF9/ABBSA9
1sQPuhyPqRFLfgP1UUprgGLust0qgbv16r2l9M1a0FSvV9f25qqLMQ3gHPTA0Z0nU0y/md/sQrsl
qZbOsy365DBuutelD6LEiS6iUC/MWeohBGofKlW/BRCe1qe+MqO/yjDfakPXHNHz9QPQ9AHPhh9w
pmT7rfxA3neudOTfggFn6Fr3K7v8QRmTK2F1e513TjyP5jRPoGYTQ/OO+eIE3Zk6/+BYpXE8zJ47
4WKWPQDvM4I/oWHA/yrC+FKltl8kJD5PGxxywPpaN8/n/ld03nU/S3K+9O5ZwDd1Ojkc8SJd28FK
NYp8fkDTuryeaD1O+72yRhENSrSVm6bDvcg+3w/ngN0woJExYw1Pwi1Pm7E018f8mWSBm5dK6i6g
orHHQLuc2R6ef7Qddpb+nG9Bi9TFFc+qHXjRT8HzFG21Mnm+BgeN7PMibd5dDE6LrJE3dHDLlGwB
PyBQHOTUkZd0kWI/si2v2bBxYx5OMQa6GhuCOHTJLnffj2rLJ57otX5hAkX5aEg2XSraM2rDj5Pr
J8y+KsMajz9moXYcL+yn0iCSMZEtQ8TK85jf0sUsnREqsl56T5iMltzb0PE3Ce3JNBTidmUyYiM5
dJiSt2+gREjvPOC6rZFZ0ovgPPAHqVDzx0yumh6NSjKiXjp7o4+zZB1UBCbsyDmRkvmmUim3GJZ0
D6BKApg8Olq63jOm+aMjIK8Aug6DvMAAw1NH9Ryiwv9+Z5J8zuuoipSESWR7aVsIBXxaJc09hBtI
/DjshBBwigpHuoR6upj26S4gyczF8coInMj17uDVkyePmYarqTyvhar5LDi38LGu032dcewff++G
AIdQiTeLfWcEIVc6iCPpdYNZiZBOmCw7Y7j943lYshD/aUBCRf9iM3WgJbxmrp1db1al3GCM/11d
ZJG8VAc2N2V0r3Gp8HuKsmOoFoC+5HRQUugBqZhaDnoDUryNybYfa5rYvzFue5mS7Kq12AapH3Le
m/eZnJcy+66jnp/6J5oMYBR/pV63AhfQoujd09EvmUDFrioaOc4gROxztHeXsXjsEo11nqdeRiWf
iN3VtIpB+vBNATNAFFeCjQ9t3F6Rut0kYEmXoTA/JUQsLFsAOArcF3A+zVAxTazkCGmnJyQ/aqiH
wfv43JDRSRTFCCp/oQv5V3x7b7j52nsKnVEluJM3oZvG0IPr/MxZrUmxj6FK8iOiTksGcrG2xid7
45GHJXq8vLpdwfdNnwRh1jbqA4vlftjmC1Nb4i+r+bULSHLefUq+96Vfw+EyrVZwFj+TKrgpKuu9
yBNaYhDXhYhH/xOFI0lQoEtjJbWNzKkI7CcDb7CN7aWQ+Ab0I9SWD4FVGxxqKWKwuCjdK7xw/YT2
Syr+6muQJjgTLOrWFl/MrvjVgI4+9eGhFhumiWJvppgfjePwh+xVHeDYg/IuFDSJuo3BCvDk/vkp
oSMOiIolV21gjPl9Tmnki+W62UuyByXgj1Yq0NP5CUZQnqbMQquO4u2tNvFZQqoPyB1RUTpu0cYt
V3Xo8tQFAJx/zwEEPQlgzTKmkTgc9kz5YtRMgfARUKCGfFzOF66J3oaFn933kaNfgjCq/Rsa71l/
yOy4Z4cS+bN56FUl13JvzbM2ckNMDWKhLPtXXO5IcgQe/xm4z//zlVZBUk/U68Y9nBCyM7nJYZ00
gAOAcYSwyB/ifXL3KixgS2J1csQxGQBGrWPXNekc5wm7vRUblerOl27CMNLBj65j6B9e42JKOdBd
yMsc2OcUoFm4xkTlFnUi48MszO+ujtwIo1A5TTIesiQn4d1qVbyq5KMQteZd4IC+uc4lfGap3Q9z
7J75ooW9qPDjvcqI7IUeKNULFnzPBDzAF8lN0hXmgBEHIAC31hQK+xrbjjRyWGGO+Y4TLk0AfvOo
+dRrySqOtioDGO0WSQPn6Um9EX0uMURAmEr3XYcetf5k+LCn6LrlHhfy5y2ck33uPE1J7++27VEi
9co78ZaD+vFNWvHB7x/C11V+7Vnv4P8J3sxPdS8wAIap27qfqp54xjNR2HxWkbPoIhwuhWJMoOsm
WF2TbgyJ7VHIGeYsGT9MmuGXx3vF5idYBLSB+jgDEjiAIBpW5eqAvij/sOqfQlTL0p2g+0mVNSBt
gzrkIOT7FqWU1cy4eFm/kMs+tYaeZaw8yeD9BsoX6oqUNL9t5H6zrwswgQDcupioeH6XY16nNxyx
dsfHeySYXvTbUTyEhfDK1MshQ+C27VOfzOAk7LjHYtCrTwZEcYknKLxTxFLfvbw37PLSQfGThO01
vga+TTMd5qfnOpPjMDmFDVLsa/ED9hzG/oKRiLc7c2OQg5Fxu96yXtSjLkgNdp3pubmK0tukDEt1
uOLkK8eLWsXUGrxYr3e281Do/Z+iQmDv84y54MewBjYJ04wDBWrVckK7wVE8XNzYvLQY+9rKkPRA
S2LSZQYcrUrfHTt1ok/YhCTVvOyfi4xw9vZhYhvSyG/eByLLYRNremtMn8zSNW+7m+C2CQ7J1eqG
rhf64M1ZHsHUvVhesJUTVnqKkx5V6TowDvLrq4S2A8cvTul5wjFH32JWuPtcsou9kTgusbA8Uc1I
Yr4//j5BI1/73/AdREsoH2ntxDlahIKvyiLqzK3O4cRHMppRE4kABl0RqqOmr7Yw2w3y5eMy1TK0
G09F1bR8VrXyeq8SfT55JwczzAAti+JzbNsJfS3Ulnf/udEe0g5GXnbsxsinl4t71Al6/5cICyDF
WyXfNPwdZtw+f2d3Bb11wejWGUnJND0utI5/WF3c+XX7czZUZx6BZescX1M4Bs2/t4iMQ/zhVPM4
n7KGciEcZ6QOCpp0WHz9bu4sAHmVi4XHZht8f8QYIaIRM/UW7BHxAGE1eG4dVWLZNzXzzsfr1jRH
ov1AGqgeoEjl1sjbLKt/EfGDC8NdKRE/G9GP1xm1etjwTzTfa98PdO9c6FUFrZQvEFFYZtsdr1w8
0QC01WLa63m5MHQ983tj88ClTq5ZYP+XgdZwOCswXiVpm8ZzsU+2thnVJnCppucQjOcWrKeJxKF9
kfzFPmxGUkUXaILkIl4/yvJKzWIGuLcf5Co3/32mpXNl9zYgefIjyyy/m3Iki25gjYL0+XIwPAnQ
iWj68goMSY1ztad2OsqWCL5KNHj3w49cMouGLLRcZF8aOumDKJgylgTj62H9/mUqN/23WpfgPScJ
Kwd/m0A8LeWqc2EY2MN4zo5ME4SeF2blQc/pn6Xd5eIhDsKPK4mB+fJ7DQu3oHaB7k2iUwaPs8N5
5fUr5DV8grsnjt/382FuaNxqsgjDw1y2ZTb6LByIW6Q0CgNpAFXfoAUczy88HB2pabPdnep/L85V
jBLymUZ3V++ahULPzf9sCWKYK1Yy8N4O6Wh/ba8ZEUJoJ7nXbCvyEq9+XPHeOdvT8mpwYJAIf7qB
1E1uwH2M3g+8VDZ5u6JmnR5VQPWpvLAV1AIFsHFGKSCbwOaBiFGCSzT19bv8JXlhjza7Rw5NiN9K
wdMB+EpzhUcE+7sJyGhxph/gSFRDnCb+4g+yTQTM9btcJ2SASZkf4jT8UmtHd/ttvco97yrQVajP
TwlozYDEkKT/Tco0KK0Fv99b43KLpPugnv227Ezw51vNy3z0aezPeZg3InSE7evMQ1O8Sv1LgXar
J/Qd+hPJFbqghcNpeCWgywaLZxsy2XfZqadGo10lnQWiIB6lI2syBZcxuqyg0vywMLl4xHYOQDM9
yoAUkaudaQansNLp2EQJppgawfS0cx6FBxjZKHYeZfblFIzaNNrGlJXnOO8T7bWq3oEJQBA4Tkz/
R4t7A5dNbHIpX895bW6/Iakx5hF4prCC74P3aFq5StxehDm3/TIOHAtSSpXWhJbGkxr19u15HD/v
0rne3Oo4fZ1j1y3XYLauvq8aZCrkjjdk2M/oP8kBh3mXO4mAsjN+b9K5LtXZXkKFNQ6Btf9VE2Ap
zx4h2Y8bloRxIOEqkA+xp8ndSO53Zvj2aM4PrGwsB5QIO2NnHWTKH5hO+tw3F3Do7WeBQDZ0t8Me
G9XVT7zoRqooc2Ppq8y3yDfhdAMIl1bP1YKjfM6HdlA97nsoYMyAJviHBw9TwylxQY6PRyB/secy
QnwFbP16vvhLV/AVdhD/ekg7iH4cah8UwnaQyB4sF6wC1RmzPXetrIFqfC2rT7qkyewCVZKo7DzB
j+YQbBp2z27D2rzY7RKEOJySTo2b1bKcU4vTPZidJbDuuyigS7JJPHLXahHpRMkxdd/TNVMlb3AQ
oIhvSVRM/ACVCE4Crm/wnh5uVfunUqEi+dEkza7rUgYqM+0UnjFhJVTAcWIoIv+2xW6EUfq1PyXg
5AX2Y9UdHy3L8IASAIQXemlZEh6TarzgwzOMZn0DGaHCRCu1mmI+D9fH9wDvVs1q11l3XYlH6lxd
N3C40tSvFsirRACH9z9YcXlXP/bwXxeppvECiEzYc3Bx3JOgr2vqMYaw5nvIQ7lUMappviJFMiJx
UVJRaT9cjoVXpDElWxmNW3eWsrqwsOFLEhR8CWZgM+kyuD/n47CM6QAq1PdkhZhQ+Tlweu8+k/bS
wAHFIl7/75iqx3584a/i+ZCw5H6Z5hdiPHzGxCtAJDE34l+anLrLw8kQ8kv5C9H8Cj5pAPzbip6i
2iv+1tDkEnSj415yBN8UBVvR+e6/m7xhTL3PSBJfHh0pKZ0fuKk0D209xRjrD4xx8a578R+s28Ri
ftP42RvzsVewj9bzK8Wy+vX9TLHiIFI+a9S9Q0PEmNNv1q2IG+v6DQfY/mtVlIle2HqduzICQSJK
zO3BeUMtY4rRTRgJ54zUn5hnqdNJRBd4nXSq+fkxehaMFED/tjJ2aFiiRceni3FZTC4NI23gytxd
pzx3hMXkQbN4ty9vn6X+CfXUdt07Pih/pcOlWNhvLMajES4ys0EY8IGkg5+p+sag4K19hq0n2YzR
gqmwsEAUEw0wYOfiulK5K0A9Bny4l7W8rsz+cyQdV8XAr9GBBt8PmMdAz6PN6lKsazMm7r41mrK6
wJfB7lf8YIAmvWkeWJ0BywXphuZhGd5VzurQLGJS0CBQl9Uq27FG4PrqkRJH9OE6ZdFxgyDQ9Fy0
+ihgfKQs8NhXVeUDpsdbWTLrDzkb0+DIDgnSY3TurK95iY5UIEpZEvhli6p6gbEIhv2jsj9rtiCR
+5Qs8pJNRVPB+eww7FzqZosZro/Qec046/5hR0CKEeeTV7ZBuwsDde/j2k8dqBoZ4T1qetvz4j5Q
Oy208yyyXn16EFoYhUKlkHAUVNkVxwI0LnKNl/sOD4XDHRn4pQYDIjFtxmWfySTI1+qS3ku12oUq
RztwgUpW7o4aaAkC+050LbL/uzEKC8ye/JshzaLvhMaYpDVFeUH8sfR8ib6haxZfc7FIcES5yQv1
jDwnfFOHJ+y32vVBVv9VsYkMP9cb7wti84M6VHwZSN8fJ62LPrzEdhcLZt5Edfv6xXBzdxn4WJ6/
jveQUxttSpJ4s42tjCIHNKCO4Qv3BJ07FlP8LscwItsS8/CVl7ggLWxiv6GthlMwEFOI1F5l5EsA
tKWgXExrcs0sT/IyvllFk+qdTM5ea9b7dWQIgjVXUC2TDcdLU92mmv9ELRPNNOBcGcdHA00bZfYG
4SGNLciZGILwUWYoLamE9pakhruXVFjbcBjTMhidHHgzvACeUfV+JnPzJbLHSDzl6iDvdBrkoErY
vqeaVa8PipexkQx7q4CCaY9tjabcTKmXk9TtFHGPqOS0ASdOqMfNU2VUt0CIgPr5v1hknB7lbIS8
1uVqVtwKWYi0Giu111/QZ8wNjtCFtYfXOA7gu/sNDSMv9I+JRTHsh4JL4b3YmyYINe6hq3yR1Wyd
YTlx/pKZOaT+R5NVF+5Q1ogJ7QSD5zx88Q+N92NEGC5h9zFGv0idFUolbT7r7j1xtBuHSayc88dV
4X1z13Otcq9Fou8bAvbCpARkwDPYD3KRUoipgdSyAbxZ6VisZAzlepp8c6HUE1RsEODcP8GqUJdO
Lzy1LEBm67LtIc0pB+uctRCpRzEO9FgHDdvEi4lDCZMbjqHKJC7P4k+dWR0MZxA18Adh8udK6pPs
n0NIkHOc/mYjx6iYoWw39R4sDDAD0+J4rQ3EXGyAFbC8cLhITe/UDU9Ff7fzCfGws9QSohalbULX
xW0niFNj4lZ7qi0Vs8zj1JQuxEoEla2UCBIgjnh9zOb3EJADpVw+MbTWA4wdFGXNul/G+FnfXM3d
SGhOfpH3OAC4nxzRmwFU12o/+hPzQGQqYUkrzoPVFgJ9SyzGZf2ZO+mFsVjmQSbTgT28qtaTh889
3TVFSMrNWLz49JDP2EJoPt+fxbeJJy3ECTLZG8N2b/PZtQP/usc5yNOY3ctdxCOJuvhSUXl1e11C
mog/oqbNgJ6Eg284XOLvpUk9uPfFfxmbMABG6TJ3jj9fFj70y2Rq0pcSPUNPTjYNj0uSznZKlpoR
iSi8bwO3wYvjlHv0xO3iCDxUi1LC+Vw7br1Paq/ShQZ2Ha3o2J9RqHsK7r3cP6zOebZzGznlLDUi
asSiIDsoLjJPXnNpUWEl8YOY+MmC40s3rf1cjbdNhnnjs/xc37HwPdi7jaHkNVrzmmZh2wGXFEZ7
vL3QXnPU74r1VNQTeBjTD4hhcFfyTdw57tKZihYRhzBdX4j6d0KmmHpDgfcoUoxeIUbWbfqj4ygs
fPFDzlDo3CIHuQMlb8DEYboUFKgJoxeDUMR0eUKJiN4YYlWlrwoyIMs2CN1FGr514Fadw5GlSIB5
84SbMBmIJNqusraHizvjzrGZog4zHJqRpFP/fnY7PeLlc6kMnpfOw7sIGi5Bw0ubRe+ORGnPDJnK
7o0jLUrxovbMfczvahW2evYsIvyd2NMGZ5hWGjtdicBCF/BdcoDg449ZRxsFmtpIKU6/WIk51Y2M
t+KQyjwH0P+CiA1kxKux3VwP+tDRqT4bi8W/RqeXbYNCSejnHkj4rsej5bM2rFuYKB0TWgMU9Qff
Widw2YPPJyodxfKdP7H9Hs61290E9ZCuQM6lwV8hu58jqOBK2PDXnlmyBfApPo6tYbNhNYErjIzI
gep7nUl5qtt067k45mTLvM266WrjhmFb2bB2Anxik2THLsxL4gyth0pmNFrU+hv+BEQ0phfk6GmS
LmFiT2EPP6iK65RRgt8dhuSoRO8rT7xdFoFvJXGWxoSMoRWQ3PNFIYe4K92CoMSLj+0wdj0CZixq
mpMG5RsatQY//1HxMj30Tfi8St9+npJP+6BSsF3f0+byEYBflgTEmD1ZL42aNg002+92nd9ihdPl
PA5pELHiVBI9Yb31yPd2nXD14a40oov6aD2y0RPjx/GFk+jf6KD4m6r1R/BPsx/8Kp181O9A3Yyg
ui+Mzeyx2SEPsMJwO5mg1OnxbSrqR+XDwVZFsbFZEhl8RBlDH0LiDGANyIi8qTq/DlA/A5gmzU2/
VZpYObUD/UhDxM1QBFPSQjyrxcg+o+RG24XE5L/Dn8wYy2F77F38cuLQB7fHI9S7ChereNwxPdyr
mKD1XBNC4YYt81xSBoxBiY0nJ11yyWDMRzz0Uzk9zkE7IL3jzpO/HPSjuSupMAFG14UTobs0Ps9X
g8Ofo/UEGyceHr1LZsoo2xQjj7Hrd/qThU/AyDN0qBDccVsthQL44KaLF10iFp1g8/oksFTggY4l
7dUBdkgY6kvMIhTOZVwMOdyhUHe0FlJELxD5yYWGJrLdE+zLWSCNte2ynvmrPgk6XNhPZY4DjaeB
Fszga/5en71LP8TdvfwM4Cv5BTTwMhA6IMZf2A++DLrqXTKRcuQOOuMck8lRhlOYlTIfEoIUzPzo
WSIpzjdbkihbeQk7zHJ0uljSCpbfvzrEXFGrV4t/LLn52M9xyIO+74wOFuWDTvq80nIG17Fb/+O3
41RsAx1Zlrg2iV9uVRz7l2+22VTa2vAFABfgzoPI6+W/VWgkoIwrd4lWBTQtewCavc4+vhDLtxPo
cHw1jUrqWP6Iaz6PiTtL42FhJZQADGtLSei/d40vkX7q5HUkHiurK/G0Sm+oHi2P5GpAQeZQFjHd
FRHxWc1xmLVMv8yd8pWkXcU4wleos5Qos3GXn0VzYzpsRnuWSBlhyugm9xO5C2wZ2ChO/B2UoZvS
ujgDYTQb9Bfz5b/Bqfqlx3x8TmeczxPMD6oLFzjw3meuUb347KdZSMxZSpVUyX6SwhUsfyeiBW2z
Xu5tHfijwUgWb1llny5zQllME3EHlp8PNGTZT9EBRyzW7FpnIvXg2KKOktAS0Byhj4WwFUxNRClv
s3xbzdiU46kPvcjWLNsfwPXAyxKFroOp2IkpqD1apjrulTfAal1Bciq7zo0agHUIi0qdSM4ihH4k
MToGWth8+ah5VwypwrSwUY+QQBZnDyLY16A1aE36gUVlUYZFgisxKva2B3nqMZNk5IZDCzLlGbpZ
X6Z8B35tYIliFCtaPxw0nFTs7l3zObIrNKLO46wEO5nukAC+tO+8r+0jh2pmQoHAjglS+ZvsT13u
PtRjtcIRpouV0hVKrhzE4pc8HcGjqQDrmV9O/rJyPYOubRBr7y96a0fH62sRej+RswxSIxqOM6ma
iCsOhB3cWjWQxNnYjuEEeJC8RrC3dOKk6M97IzW58mHU+G1h41F6eNNC9ohHcGIgnzkhcmGUgW1U
0LCFYJAV1DDq3y3/j44exivl1pE0ItQfTij8eZDzIaurE6XdQkPMNTZcQ8MQltlezT10J90OWZXA
w26pgMOtjrdcqgfxw3aaNXUtou3M47a/l4nbL5MozOrhsPM7uhoPTi2zn5dtfr/FHTU+wFxaXgEW
J96OmG+cWfmQrw5VjrhVmzuHc3GF58MunDSwrAVgAyPEZjUaG+wjuS9hrp9yb+4gQk61ZmNtRAhB
FEGB8Op6DtPP3A7jKw1BSxl9sR368D+k06zBXNg5FCWOK886R++LfWTeQG6MAF+H29Q0cF/AUhVn
w8/0WMxGvHFSkxDzJuKZroPezgpIMQdAwWjSFVcuZlglbHlLZ9DDaVTFOsmokN19FgxvGpjOXLCw
5Bb4djw0uQkyNrWuagiF6H5JYLZQyyNXyeMNA2JOWoUXqQyvOcukngxKBHJJgFy5VaE6Kwjn2PPF
qRrV7UiQ9N07ADVncNNGHlAc0zJgqdQHausda1WYpY/9mG2y20IIk6dePoLcBTJ22RxRoitxna4I
nfoe/Hkkz9+QRJ75T3o/BybDAQxzj1WgtyIN7DRE7Tdg6b5R+tITXx0pU0wOfHrtO8pLlzz4VAFX
ODHoIroOCiHC99VPZc5huBN8Lcdrp68YZZoyADU0zs7sQXw/NTS+i1W4wJDTJXe1r9bvAtXqjZZK
hj/pzdPUNLzvxS1+yO+yh/7fcnWi9ET4g3jppRHAR83OgpLGYQljiB8wb/Cr5Ajpei4U01bk7F/c
2JX2YWMWfazNeYwNUFmjqBkD/o6qNXfKbhiYG9OnZ3Vm3b8KPJenxzwd/z5vRBEqmLWKRBgOevN4
yJWKc8i4iBwxN6f/3FwTc91LdPfz7Pj66LBO6xNWgZWCLF8iCgJUH+1cGeRL7wJLCoBa4HEncWNO
qiI0ssUXRT5KXvHvXlNKuVVwS3+5R3uKrJ3WhvblnzAt+kQSOacyB95UKpKhM4z1zEt3RMEQIJMo
J1ERASGiuLcgu6PfqGNQ4ekdf6IOKjgDwkH2mSrAm2IbSr1sVCqzvkgagg695RRcLjJreC3QVjJ0
M7xesOvQMMqeHgFv0gGX6Z0LNTfouVrpLAe4IB9n6wJNMe7q/aUTOWKYExHBviI/9N6+eASRJbTZ
A+imHSpNZA+xHcEuA9mmXVzxVK0AKwEroc6kzyVMy7g2Ep0v97+RWUUE1+wlHZHIvhng3w57XsJZ
bDWPAI5h3n6Tcm754CUThY1q1OuSAU0NpgN7eZQoq/W/GEi3dWgL8Q5f+b6oubAyglcoGnJ5Kpij
tH4qDTlwpyew/Tb5N7vqClJSNmA1lOcd6H0LWsImH31hLLCavC1A+0R03tGZJDP7RCAr4+cg3VjM
fJuyH2CvYqtHVyQ6VIo1dm5nksNmY11HENedjI3m2yS2nE5BEevgsi0DHs3nKLSfANK5ibIjbJUv
dFpHnHtw1jRLUKWrTWgy5pes3zvt7P+Ulx89fobtTxuBuBFAYs18ZyCeHvLKN9Jp/1EyYI9o1B4d
sB5kY33RSQBd3mY7iMBfkN/iFmyBx0I6hz6CcCY4kzY+5N7wLz8BkW8AqFsQWs8uDHbiYsTXGJro
+lxZ5tQK+M/rZtGslz7o4G0p1BUZokCHJ67KCmVp3Q6+JHvnOdANqaWzEUvLxfVInzpXILN03Syf
IOKf5+ZnuCjtlQ1Uhv7LHyk7J38Y/iIsXrM3srLwYwpGUAwWk7nMqfx5lhekaruuL9TfvDHjIWuc
qYDutT/TefidB3c/9TvzWjZoccGJB3gu/1g4WvpIrEyy8iR29B3ZQPFXnQVKowb7CudjiSiHdSQh
l04QeLs1mHqe5/GiWG2OSDPzHyFHJe9pVpXKXRiQmtHiobTfRJytrfzIE2nJ+xDWfu/jRaPu8386
VPg2r6YbLRXsKFn76Xbn0tmDG5goTK8ggJbRK0YApAe//jZZ7QjXH63rYItmNTsxcjSrIm0noHPu
bpZTufR+XulXT7V81waNwyvLXftHcIbXgPNL/RE8qUwgzIfsSal9nXCf7MReHgNCb5zqSWbJqzjR
socEojjULNHDh47CuW/WWdoJzmgrZXRYIdzWlDbfbO67GSGw7uJLWx1U9tsnHnmPDqvy4Omfx+/M
IyeZQcvMQPlYNppU3hiQnCtUKCExeZoR/ZruUIwZlvJ+uVqCeW1hQZfU43+OYGrZeYW3+oA44X5Z
frOlrzJAbebHt7fpssY8wtUsSrRHGoZ3b75BdPh/WkHqPrJtNvuRND2ahbNWUF9frG109pWcb/Lo
FiUn/9xFIRQuYa8vLQzbusl+wCXMaBYJLGuT4WiXIw5s+wuPEeSTidb1s4CZiPqtu8M4qNgIjOzc
oRsn2HsEYRC/QqV3JSOsnsrFSQeI4cvDDWlx0pPeh+JC0e/WfzaK5i5BDzoe2zrbpI8u1chb/Xed
jPSa5bO02QET5d5WUxZ3PQmBweiVgwvuFfVI7A3zWYp9qrsNxDkNFFpbKVgZDbkjejtsFVu/h9cB
2H+RgwDw6G2NUXwz7QI94XiGzUU6MafsNqYLzUuFVUr7REyFW4QC399Bhq+gS1d37p7ZlqLdygzy
duPbR2nQsaLGNGWpaLvWpZ+SJcgQRP2bdGl/OixQG9fFl3iUVUD2/buSAukP25C0b6jwppMlvPok
Ga8mJxyAMSWKI05WTXfL9MfDpMeDfGY2IzUxYH/fTlTI+r31+Z8iBEIcFVVAMfiAimpJyAoYk4Pf
bRvr4DYP/D4cVm7/DGe+BYdAbm+z/V0xuIBgWlakM22j+O170BdcCTDqrDfz22i/e8eSauQo2h/S
6lk5KisDvtR09zEt6+0jXROyd/cgMlyMhWKvuKdMTh3dSX7rM+0yd3xZQHzfULpn4r7oohrAZoJM
zhZNZtUpaBZtfg2Wp6uQbYAP/LsGbjcXkSLKy4YIxlIgIe1O1VF/suvxzKxgWuf8f1cw/FurzDwy
rVXRFqtAmHdbdYY9IF8mno3v8kt/eGMnxiFYvh4DlufQaN0WDMCMf9IUyJuUjw/dOquXV/ubwOwT
4sO8BQVu0x7U4OeHqOywFrxNiGc/7RULW8hve/lkxNnuixxYznxRQMVHYNQfs8am6mx/Smp5J79x
0gv5iOUxCGNmtWybpLeSfDa85peebcN0xDwORgqLgdsRexG3Pyyq5Pi1rHW3TKhdXXshQE+/FL9b
1OPtghO3Jwo03xwbuRiOWUl2tCasJCrgZBKozVNHJHGxg7LePeN3WUrvO0oBSMC7JEaNF1Oddzur
hIAE9KKRFcQTUOFUVmnKSBSScbka1JgVj87reISGfxUHkN3zhgRA3387fFO9TvBFqN8kgpx8NhJc
LHA/n3JYZk+5Gy9U+L3DBtvQTRS66ryzD5ioyZ1IZ+7gsf25PoiYSZ4+2GoINxGnqSrRwWDcPHn9
cHN2DbPN26Cqda7QUdQnlks0rRwNhDPCxZKh3ZjggKXuM1oExj5V8nzh9vHu7axT7UQut4zS5LE/
ULRYzWMf1sI29HKiMBjbo1LkYM9eIwU82OST6FlcnxnW8UPuqk1Lj2+xg2kzDH3UIgCj229bLh9X
hfTtt4uVC9ASW8hl2P+sXslntoK/t3K69SkKg2a+W/FmHigdt7w/9Og3rdtdwfCOInyojBZGsfbs
mFrTkHa9hfZoQXo4/UREE1mxi7HgUsOegGqfDjOjhXTp4RbKnGhaCZutUleOzRxgvszDQhgt1bhT
byJHT9v3VVvkz0qSnAdFBGTQ64loFFR2YCqOQGl6Q+P5xellmBEk5yR6FOt0kuAn2HSadTpcBjmu
OFt4IAKHKHl9xsI/WTJ4kq/Na0ACmcfBGAFkDB2doAY4yLYqzrmjgKzb0LVdLvEWlpLIXgNIb8RG
Keuhmgdrqhe/GjWTIbCZPVA+PNOYvDhkeUQvPdYkFFe/Behm5MpBtvBTiwePbYAgNl3MTi7LJMU8
e7YGv5l4kEbnkUv8QXpFKRV+C1LE4OfUmjqGTUEnkJMBqBDWIfLtmw4PEFzoz1kbA5Yn3guhbPOC
CWTEFA+n58Fngqis8IVg2WpFT07/DVZBokj1Z7X6o0ceDbB2CK3Cj02DrLF+DcRa9WLmrKEa79UH
NH6hfgo+tE5Nd2AWQ/o9oFokE3vZ0d6BajhW0HWMml0tM8G4FCSsm4zHAGmjDpXBQuH31TggJ5Dr
k9WrjDpUS9RQFP8fzvomioNmd0muiiQQvgdGeUZwAYm+ViA3S6k3BerH3GUwe95HIn+3TI0k4pL9
sRF2Gk1r/9WPBlGiEkQS6W7Iw0RADIWDUW6yd7SR3IfBmpWpiQ/VEX7qQSqkO4aTwvNpWoCSEXFt
Z3YuW0nVjBTq8iLTyFbdBWu6K45ONm8t2OF+itPY+gPgLP70n06q0BEdQEpGZX7W+h7/fPmgYAzV
Ux2TeCOXKDM+2Rwc8u8O9ImwDTtrAlnvojAvchedTvzHdQo0GJsSn46iScanQrlg1cYuPJo4h8HV
wTGbhFkKSMiJ77VxmNr8w4khzQ7maVK+etyMgLwyco9L727twCvsaxEK6iYLcwy9si8a3KazuWK2
Z06qtmTekKAedkBwvVBUzaHBRMxI4+bIseVXtWcE+BkIB4N1K3xcXvCGME4OVds3TrTB2mHwwnl1
7dUIJq6P3QdA6zwUTeccRRP9/HARa4mE26S+U9ID8N025W0au1htgLHB2r2Pv+F0JrIJ+bJdJFSr
ppSvTWDj7jO8+0CydNHREEvWAMm1QdyqJh/RnlvhYOqhnTzd4cQOqaVSKF63saH4KXXVRWJZhmKB
JKA8svkydu4Il/PKiO/wFceysWKHmBhjj2+E0ueSCgb+qpcG8d8vrhMDOMJj+p5ypYgS9iiqpE2G
97mlDafPYu/ojM1umgPT+5Gkm4cFHjQCcwc0Wa1oPqlUrL2uoVlnrCkLmBNew9QCTTE8KA7YPnZN
zhOzmYHzUuf/lVjGkzroMyi+A4aN4ItrZUZiRzDxwBA/+QNOZUjaYv+zARUdzczAth8iqV32KAKT
t1QDlM5usOzkiuvnENKBLPN/H+mgHTDounUdpbzcRa9WQ7i32uWbDL0MzR+Tw0KPnynvosSBIc5y
/Gtn6O2jC4Jp/56VoUOiD89KHY/+8hcGnS8z39/+v3TDms9z2oVGEKhALW/al1ahnRDL7d+lVGxP
VI1xk0JLYEgmuRMd3cZy66mXleqlFpvDmAf9xbCapud/9/EtXwctpjDD92GtHYbd9SX/TY3npOMu
7OFCAdZLjk1S/zf0kIZUpEfYpfY9da62Mjn8J0kBRWPxNuiQQMUdLVQ3pgyN2/cO+uKleOBJuANi
dYjLlogEOE5bkFEFMSksbsvmS7lD3addDRSm83kYWwVJ2bCe9gi11Nm71bHixpFP8VL0dZOG2gXm
S9TKgA6RSU2jenrlsc2ULuda36fcofhPWMw633Fy0Iq1TfahTm7/M+1456LNCdeXS1iPB28Esw0k
RVFNftHsv1PWnFR+i6loud53ryonPIGhYIF0ETrPvglk/XR0xSZ7PifDcYwVy+28wM+vFwYMJzgD
qHTaubhtR1k6i9AKgk3m7A+QVrwrVaveDmZt8zzTdkLKPoj7W+y2QOAmz+mLkNK6CotN2tPHe30D
9mLP+WUcEDGOl9KRYQ63jIwsJwDhVRZL6X9zKElx8R3TV3CIQe7qg2MVBXQrK9pWvkslJgHlyJ74
qRz+hIyWz1ejTuwFqK1Zrvtr6aHFUcHUgJQzRww+yEj75iC/oCvEfY+PB1lbIzaAX6wk6fuJthyE
JdM5FPVKYRlVSX5B39BpBqQuI5pEwFDN06jc1IwVaTZdWuDFFkA48DXHQHhuwXZmMFSM02BRF4UC
XY30pLXQiSx/OqfRBmAbuqIFKQNkwU4LxbhtuHGo2yaBtCGdw1oTbUOo4bO3KqhximttbD4Ot7l0
zWiviH5QMykE1HeNBZi3QBADTZGllqYnH13UY9jKhxkGlxAXY/9zCrnY8VVd1o5RZikaKKpGj5pF
D4k3ZdJDgyZfeJq2Nh81gdn/GCFhxWcJc3lcNlhVxVZExhXL3FqPlL95l9Bc1626KQ76bAriwz+C
MDWgLslE+tTIrcCb4ZiSHHxHtFvpTLJzsNsR/KTndPv0qyFPptfDl4Igc2fYHhQVGYiDVceqhgYf
yxCYPSkBCRNonuytbw1MC8f2MsKYaNlXIGcwk8blENeL/oV+qUBireOss5OurQtB56qHuu7jbubB
xkzrJ+J1EvZC7NLQtQM5dZanoHRxgnoTwdRqaw48S3yZtjSynRHlSCitcV9GbA76IoOINmmrkbK6
ZIpPVWHQbhbDX1oNZiz2Ygq3nGQdxvg+pE0CLWyYvbcJW5c7dXj7QvOIrOD5uaAGu9+C8cZHCtMU
CL5nCAOVmCCfzBJjx0UrSihnum/xSZX9VnoLJ2aV74RaudICcKOxeS5e/l9heaMUbBqz6JQdzxws
fdstwyyovA2Tb9DqjWUoE1wFMbU6Qp0WO9jR3zQBwL68q3wp6ei1ZjS7+3AQmEZj4d6mRXDDY/PD
PhuNvNifRdQ6eTV/2Sl2XPEHGhSDlBsDMaY1tb3Mjf0KqdnaftBW6l/FnURPMEAEQhizuP0hd6Fi
lw6AIKNF7ylnB44Kav7/E4cSxVtcCfa2Lpp2CCV3utOKNofJIXqVpfPWwpib7lgX93uuR35mtmDV
OCmltVDxL+b4WQBlnR6p0OckBVBtdFxpJxj4DQM+/jvs454dljG94vfe06t+kUTEy8/ayaPBul+f
HGMWFjY6ZRH8/aYZG9w+6urNmyCErh6xbjiwh1Ig0kOYQBnElZXJLNfWoIHKs1NkuqM5moc5Ajfw
7sdDbzjlTG4n8Ozo0XgKKLUV8GD6DZOj0w5gAlwPdNmLTpjkzj30ZXY9i0QYWHWdCUWrGfJiSs+/
qNLrSSPl9IPNnlx5tAlLUlv1VS3bclW4vnxcAcIQSSdarncTDHFT6AwiilMacQkr3nnkTYXOEga2
KKas+SjcWeFkmwMMaT6RvMP4cgDeoEF7OKzS8FdieaXAKvacn5c6dhxCOVEZ/1vhT4GFG9y1vFUy
93VIjGHYyKyDgsj243MORGQ7VyQXWkCmMFhjLOcti9rSzcKbLAnG0FSFC2kuWtohKJwEAeSOGJyJ
FiVPXsOiABvFcPn7y5j2dGaywYKPddvS1goB4ma0ZhAFrggsqPIWF7mlFxv2jyW1s11VSuu4vT/h
W6C3uGr5c0sMrI4SzMB9GN4Vauv/bVzxFOYjl2HCyStvxHdkVZxRP8UTn0bogMlnDQcEUZhs5+Wy
C01Cg6+l0X5W84z6nZ9UO6NG7g2wq5McA1wq2sMR7IosahG8/3AlEBzDBIrCc1FKp951wsHoKxiu
jOfJCZh7TSZTjfLoOLZ7xBlzDuijZ34jWiQ3wUTR1SOtQHn68xGY6xfEUFjKtCx0V7QmkRQKTVhO
n7wXEbFm0qtb7ZZkqgMOhBCgwbj2rUgJYlAG0Vn4Cr5mWgGpzMGcMy9wZbae/Un+CFbOidtSHo8r
LqkkPfi/cvdUM+fRYChBtkxwMGubM6t22MeO9kMLixPbIjhkvZAUOdVAQP2xsmirpznO84NVIHYN
mtVs/YL4Ep54oj/4YT9JioOapLjUbMyKNYD1F4+cpaDfDRGtARGMMOkVazdHOdLNH+dyokc4ZFl8
Q25sscsgJDAdfi1NS0H/xM0ScjuLdFIjq+v+MQyJi7L4mhDwHNACaAVyOjkjqJ1O0xrRHXjS7CKT
1EAPf0o2/nliOIys0nOq8ot44ThWdHmd4EICtqqT9nI7ykeEP/FLAvu+XxDCv8HFsIvv8zEKBb8C
BNZl1LQrRdCu89PwMulcgga436N/SpLm173HJgceDFkVxOveaUUjJrsocnfrh9D1VeFU11jLWDuZ
hrCDNVJNhN4h8iJpcMLnGsCYaR+h1Sy2oZSdZ2iUsZej8AkNFISuqMrQ1Y53j3UOF7M+eWnaCxeh
bsmn95lX4Z6BQoj255Doa8+Wxbbt0ttq8EORaJuPAP5dMBM8LqART9u3lSB+wDAGepVZIxycpfS0
o6Uv2sdgIiaFdOMH66BLIkSaqUW40mQFoaSNibJnSYDBwH5hAs4aumLRM2SAUUpLAQSw5bGIxVB7
SgQ3Bj/Cx+bNSbR/zgSVBNAqgrCiHVwM4m7mYLBOonl45IotocIXCSLlP6ynuGrqNeprIK9WF6NW
p1fM21tpulMVw5tptoydGH960CsNrrOzCvKUlvGg21RKh6yMlMWNUGXG5QzO/tSNEIutHwzIze9O
t0lnd2eWySxBD7pz4N+KIgrJCE6Gc35KBy8RUTx/H92VEIQI25Z+8wtT/OYxmDvmhBPBnwCQ141L
REMBpRB9niTptuozVZuhawyISwGn5IUVTWADZn48FKa5yZkxcxtDgRTNFev3bsUqID63CIHFPvSL
A2T8ARpHitprkQXWhw9DEiVHeRHXqWVK3/T/JiqLxuKoHNxNmfdXLbA9xPIJWPkepXc5E+t8H/cy
Gns102u2j9y72oFG6LZcz7DIAorTY3V5LjX96WHd74zt3ueynvisVEc8qIJiCKWxqcEb7JA5q225
F30R+sMxhFksPSSeF0aNtHg8RDOnhpvesqiw54w/2Td6uZk7SJSPRuG6uj1sDjzLs9Vdw1T0yAgP
Nd7Ymm/rer1zrB20IV02SrLnZbdzkrum5xBowSEVzyc4X6gHOf30LvAE56d/4jQSLPyzmRvdNdoB
qphaFDIAHyhSIPJdTV7pINhzs9y4x0I9mKb3liEkJ2b4GtAyUH6kjFtvMQuxRrlU4d9Cc6Z5rWH7
Rwok9JJcBjiaBXbYQ6tfBEpV0in95noRtI/B1GXmXk3F+FH7I40vBkK4swst9PASm/R2XGQ5iQ+0
B3KTFO/CiP+aycGBaYSdRQwcnVMxoxwAzohqbEjtD2OF7aYve/+ouSYMDR423XcnJlYpt0mb1K/g
0F7jlU1HxRriyyNx+E/v+BczxygpaTzNW+GMthX+C8nO7Pp3DeRwQVMeBH2m2zq2gsaNGkWPVBGV
JX/E1fV/SvCfF2MM3ljnC8Bk0H2S+tCgYrCz+22vuxAVDCCGhjKSQ5tW0dPydRMV9lTknW2FhbiC
CG1nZDFYz3NWyA2/3+IQgD+W02D9q2DwAuj15nOeG+6N9w/VZZX1C0akPEyuF4HA1WpvIbvHMuMF
i50rOLhTrYtZIrzxSYiScWUedx96iDny5gy5QoemTuo0RiJSjsMUHuNUnzMO1WyuIty5TDbsFtD0
BfR/wLuOdT5LRqt5NaQGREgSCaF1A2FPbQXG7fjm+2od6K+ARaVpFRZm7c5CV2sA29XKxmyfVifK
KAHmUO0yzpjyNpflYUG8+JDdPDaw0Lza06PcDQDDccOEYdE8XKNBhC4Qb8HNUkIpCdle834cTHjU
JxYTHO2UvSoAkb4gutvkn6ko7a+z0lCZkTiDrFyNxs3dB6rK9fYPts7iC8+5jG8c48DyEnuC3Kcp
+mXzHQTo6I2lbJgHJM5PU3N5aNVOE6ECBaeITwsebHoHxPu+cH5KlYv+10FRw+KXHj4UWgmc4ozF
fwKjhIsKSELZTAmeOJ7YrmaSuKbamLqjBCODoGhwLfk7uzC2gBCmqrFAcsbUwwl3OBMdQhtdGyBM
8wJgKWID+IjqBOuEHy/nsoRtR+ClPzUZq+Y0Eqaa6mHyMw9uFI1VWbYK7e1Ob2lmYOEIi+zIj51Q
h3wEEGeclTst3MDCzjtODEwrKA+D67GzWEv/bR39/L8+lMwkIHwH8+ewL+nhUVV6NcYTGtsxokY8
FZfW4sW5i71hl8IuhjGr+4URH+ATlkjthl6V//esVm4xg6TPBwTOP1tqzllvXu026NvmQS3+qqLE
j6aLI4Tiy7Acf3361oRpbc1c9qmHsGqUIBpdManrvVHSTD5fqPb2UMHi0hGV7TWGRH82HF2bnZ6j
XNzNkHnele7UPuReDA96+OD+lpgny81Su8giFe5w0qkr2CZjydHFFt3VMeJpwCGfAv681KobdJKN
XQN6KdmZc446sLdt3Cyh4MLEunHvEpI62EUUMitwhDYxAqwWCui9Fl7Z7Whq+tfOuv/aPONrHIFP
wT0fCYaDe3lEpOeqIFVng84bDq4aeAKTNkAKmhrHw2hwJNes/StORm8XebrykQZF4H8gqPxLgiMT
xinSo5bORb8jIwX7tI+YOS5eWMaN44VYfuo+WnPelg5sneqc9F95sWUIH1/ZCcIhjpHe2mo1YezT
rFna0AbJdZ5lToinsJasSs1Wz9W77VA5jzuryAPBiJzm7gBRZ4cNwrChCpH9/Z7RKVDAtnJ9pMXf
5JmBUuCz0Qi4t2otMWfwMQS08fqRB7ZcsNmUPHWWgRd/KNMg9tQhqdUxVZVcHYAJFl5rYg7uj6oT
7waceyuHlE8ganLAtR5tKn8qiiaaBNhAVkDDClVS/fF7ZImd2ItbPqqfgn7LuDSZGFAA4L2HyurI
jNBXPdlwIWVmKaiY9pQwBMoU2Lv2+4uy7huI8x2Wk7vmAw71LCOQGjr2vFpZlz3CYvXLS57xUAv2
/TPABmwjaA/bRBoHLCKKZo5FKdHz0NVXMRRbgk64ud2Lh4PtaVvA/oC3y99rNHkqD4T9IfulJBEv
apqMratAUO0wNWD8PTokj4YQnaf0C0qvQWBtvlx9hVMe3O/a9RFUXtwkX4lVp2y6hN/PXY+oP0jv
WwSegmKPLfg8duuLZWQvHHJnlUsuZ+807BGBOuIBOImSpvxBeAi3rWML2LVs1kL1nOuIrdKQ78FF
SYAg10mdUoFtYEetdEArTuW06xy+AKJkSgT9iduH1EuWyLM0Ykm3Zs/N4bRcG9CeCWm/B01ywY47
yS3G0q4j4ppV+0IaKVCEhpuMgoLwB5up3oAfoJai0dAL82Ogqy713F5IHarfW1tBpDFLlNDeIh31
6tWHT/qKMpOmqBVo2l0embKdUG8eCvQdQOVbA/7oROVA+XcBL8hFdN6Vw7cqkSmYSW07aedadDWD
SP9o2IiaAncMSJDLAkHxvZuXR5SMuFIIClYraK8DdqUrrB5CHnj/cihrT9ppPVnq7J+r916E+vF/
jYs2LTHdAQe2KqG28DXRwu99Iw5ZkEHdIgoqhmVJ+j8sOOEskqhVUNOxOZCKaPm4DV0LJCPw5HS1
1Xj7pl49yYnSqsuzNiislLDG4LzOHi/gO9Nr/YzC8cTtHj5Aw8taDfqHW+29Sr5gqeMJVqAmMOZE
xE218x3LKNZOsAJcHPv+Qth70+JR+IrzZLXOLXfRAoB/D+dvJQA07Ur3wW/oS1rAwkaJ0cvffup9
DOy6dVwJeyaiZpodorTimQCL+9lXX15MDDgo/diDUTM53bnjP2c4Ki3LW9d1eFllDH6OwC+Zli/0
FVtqWTIAo04yCoIStxp7CH6OCweCE/lXdxx4UBoVSWlS/x6TfZGPff9YHBVanNeUyyWrozcybHtK
qmEo5mAELJMvgjNSFBmoQDuLBnpvE3zozHfCnYpWtOmAluRV0IVNcXZVIdROUj72mN1RvlwaxaOk
qoNXppz7up/VzwCN+PJ68cl3RzGFH/kdaBo4miRAVnpfN/duqtnNRGo4XBp6JnXNjse+RSFlBlQl
W4dkP1QKiOibEganOdzvNMTjffEU59FeymJUxEciFDf0ezpKFHc1u6LadBnOx2UVcklKNMzwtXrB
GFvoPzgr0zOxxPMGMQ0mFoxkc8vLwCqqdwjtpGCJF8Q/KLfc5xZPpWV6GhIx9zNQ8xfmIlK2GNll
2RsjglxN4zLvvFFWGW7wdDBbVnl0/JswYcLqf4IhqI0NV2VQLvxF4ILvRbJcNeTxV7OwMnHnbqsG
vPTVdJZekHP/9dvgkz0kElcpB20sSTrlbx4dlEwwtGbbC27G84i20cxquJxOO6TyhvLu1ymBAzx0
aj+E2wqfz68ZYDVZlbRfWjogDB3UXsqAd7638Wx1skW8WAchU2n4bdnLE5+M6GFI830HlCMaDXmL
7VVircjcup2QExyb3OpHCatdl8Ey8aH+Y/qvestYYTROVeAX4t+mY45/mqzt9q5usux2J/Q53zlI
G7DGzWA/8BzMpZBjthwhf4SVrDtlOGePTTXeoYEBJ7mqqEvfheWOpb1GuXGjMpa8pWmvvFUWcpH2
De80p1Ff/9yBF3G1bc7lDJYMzBNeI86uvmfE7VsnsZUZWimB+rOY1vYCy169KoTQ94P8wg8uhG5f
KWMSSUaAjFB0OZx/tbtMk8zj/1rT/Z4oLBSv+toPi25k7OqkQYXhdaezKlEFZ14GROb+CMwnGwx5
6ep319l2nPfjTmuSK5r4Ly7ogln7mBJoImt6EQCGkq7vdwKlW5a2I/uSszwLWSiTfL+iGSgFEzFJ
Npddff3+LmJbVBiFzAvil7fdZiYGmgM53Fm7DzgE3qtjCwALBnNVNSPvnMLidqDnqoNhKDsy4mIp
4F8wA/61ORR8vZPUaOPdZM7LptnWWoNwfIfnY5rgK21vdJdKXvWHs9OHudL5xEaNcK5KI/Y1yReC
VlHM1roqKz1wQ1D1WOo7jwO7xu3hlWGEfh4s1GKi7+Ij4vAGJBPbRviBc1LVA6EVV7HF92i5CdPJ
FlNv66Pz0fXZDWwIAlUQG4DVMR0Jfga46J2eo0rop/sNnGi2q/OjM+4WsU4vZjeUGrKuqN46BflV
EnhLurWvVK5YYJzB2JWKhGfCCOXCNN1WVj4hOiSNPu7hmeykcZn5cnhoMZCVlIVZofIVxlVflT59
ZB2mrwaUMM0JLiMwhvtRNmPrXTs3t8q8aiPp6uUba/fo8jVaI4W66oWqdXF//5An3h6FpkfgVe7i
3nhuxEWS30h8Oiauxm6rKKyZy/BrF+R9lQ2ShcO2MRgU2B1wqmaSsRFNcCYql56zjQkrLkvLG52M
NwYGbws0z7yV/rlqdRWPYcXS0ElTtDe6U6RfbX5cy1VimQDmJWiYUc0G6eoeFk8mkbAs/g3N3Nc7
r2PFbZNPzqR5I/7z+JNHwz41ONQZa4gCVswzJpF7hQeECncnzxe+SLOaNGCCX2BaRmY0A1pKQ3YP
PL3ySgWilQb6zDJgt3LhYMI0oaBkMel/LLQJG0HKFzwUU3eYqxE86PIwc1Wq3tp8bA/SRMiXORUQ
BGPZeR96tm8tc/MHJYHQsT0GXp57yTxocuugpcyCAKApQ2fzmrAXPDq93EM/5nFu3W8bOZPRbKSe
t3RB7I/QL4dx2PEzDT09vFM8nVxr16mm1imBCFi/+6TL5sG7jCMH4vrk6XYuhXECJQ78OB99bAvR
eAB1gh25IBytjR9wEFexLbR3o92D9r5LlWnYY2tTMS2BGOS7sR0Qil8e37N4J6ydxe7rkvm9Ad6b
/HS0HwhT/8XFqY3n3/LAtzqWcZ2Fcsw2UzTjHPxr0MGOYtNnJWGMBcZXXB1DLhooWwP7+uPzhMBL
iy/BanwHiG8L0gP7y+Vkp+S3OLZs8/iSQCIl6dki5/zEk2NCxADpA3AlARM9NPfcsyWTTtYheAVB
OwIiLHaHkgyTKmMtjrFY/qJC02d7hkXL8IiwipBqMaffeX2JjPHcoyuO9TPSS0mhxAuzPbcKDIRi
hcTh5GKO52CPAhCDM7liBXX7VjMODvhIVfSHSe4Om99JTRxZvH+NBWiDZ0+IS/+gAplAJCCKydC5
TRVVqH7MrWsyN0lrivw8gE+Jj7uI9S+DjhmognXab55TU3hHOnA5xqKymmSP6E/kdG8hWLxaAjNt
uWkK7T3zLqLEK1MRm565VZwqeoH+AI3ktowItg1B0ntIKRUdzS5N+0FlEmR6frwfa4CmarALu+6e
g2YHCUqAm3dtsXXGIOUzag518vpAIJvLVvXylQTLX4UswMKeNnS58Fzx21rRN77RTV3CWB6DM5/y
p+JH7VrOebVt+uiXoGJs2YG1X3cPNurv6WGKflhq8c+9/K0CuUoY3swn1lMBzHg2UYQrat7YsrMd
9cxU13GdQACWYYEZz/6OT4C/E4m5CMPp0/85M0sYSb/QZRCm5BAG64IY/UUBVJj6AFcj3xevgAZr
+2jIOZAbMyeIVFR8fHNYRL1rp8fM3IwV44NSSD505zogKEgdT3ktIf1y+EV2YS9hQdReZ3v5UFMx
icYx1GjwwHoc84BpxtP/PEnl7kLCu/cDqEifeahg5uK6tf6icUErRrATHQkmLB8w9Y4TjrlPc2ly
UZ+U7KG1em3lFF8/E9U+PMtCrRwy2Ygz9YLhzJ7fTrMK0H90g7PWJebAhSIEHqxfna+p1X7B2sZH
bYZw1f2qINRHW39UjqQlF8UZMV1VKwQZRfg13u5R3OFDzOcxdu2s+6KwZjCQZMSn9Z8EG+LenFV7
pC8tvHtEuaSDwPQ4Hh1ET4wA/9S+XefEt0emwGG3PCES9pzjjPG6OXZjX3geJNmvEr5H/Pusksqe
1KTli7qfVGJLLaACsf5qYb7pb/VKNRNddqJAHzNfabX5CgFo9NqNCQYkweFQpxf3pnRxOjByrMno
datNWiqCgWOXVB/lEDjlqzWhHALc6KinXFX9n4zUDMNnhUdJRfosMvpyZa4N/8ARaz4MzroWmS8v
sOY7Bq+6HFzYhcg3goZP04fe912N8QFtX4wOzwb2IB9DEwMFEqwO7hVAVZYS3Nnw6YHxAwXgbQgm
honvhbEx7Z0oPc0+l+ItcxunrXch5IXkSmUwBLwqJlExk5uL/wIGuua+EB8Ad2UWnnMVuaMKDfHQ
kqQyXk58tm4lEdWsundPAhMqevEpRElGK27qWGxv2QsjqvZJl9gnktNz7JaYnomtQ8WMCvXGK1qy
Aq2vF1RvcKDV0fEgRs1v/AkBPcEoC8FkdnPlTEcVjVmHuFtRnkTKaI7CBSqpEKcysXNuO0hNinJ1
KevRm5dknQ6/16ateP1V9f+SGp9eTu+l5cphVHSluK93LzzV79WbvKQOeKMYC7ShvgVZGFb1rgKI
4dTboAOTFigZneVM5rx8MWeoBlv5OJCU3QCOdhF1KfPcNKPJDlH8p3rVgjqobpx1hJwGcTEisEbw
lPWkrtDpsEGLCpxUthC4pM7JkpZxVvupmOZ1P14mdltDLl10D3Oyu82kQ25VXipHT35EtuvVhrIz
S9n53RugkbwlPz+Hqc/PcTpn1Hid8FLXdWGuvCNRe5Sf4WVozqAFztRWoTREwfO+vaeUcFdMLYH2
Pic/WCe0+WhDe6E64ZohMk1oIuDkyLBbDjThLPX0Qx97QKc7BAdlM6agP9fX3WL+QF/B7JM3AvXX
iTT510HTGs42YOrWIeZ7xUesbNwt1lwDQD1XwEEYaqhvmOh9qu9Oyd4WE3U207+woFIsZG8TJVq+
pTQR3D6Epx9eiAJYZ/xBsD+ES9hH4ZdK0vtQQRpKF9MocrNPoJD44SAqcIBoXQvQC+zhwo8TJXzy
/EmKztQgKWNzgvk01GxaHvnKzJb4fEx1RdmTgbsZy5SeXGrklo9SNBWd/Nx7UDCi3nWct5cRjlMW
AyiViV5NUQtu/CXgQC6ACqfXKrL7QE49br9gCnCK7Vb8JF0HRezeYSR0MW9jwS2Q629N6nMqFSfe
DQlOG+t2f6iAm8cUnRNbxYh9zvTxmcJlhTq1A6SaoV7taAH4D5LDhYSRjnKnOb1RILerluwpL6Vo
oJ0qofF+Lkq842e1fF+7+odS+sNr9yTrVysKXsPgccy4w7x+xEQoK2/razmIhbhTlPIMeP/gSylG
EUppOLHwpOyeAe7+N6GaiO9Xjz0ly1DUuispe4nELqN4IgdIYg/p2o0o37nngT1yseYg9q9GVgFQ
MzLX2QiULDM75gkBrz/YQ9ThEt53f5nbTPDqLokvvpCp7SZ3YdpOKWCgixJUc7zxDo6BBeW55IxS
CWDX0DBC7G6axoiskGtoO4SlxMYX8zoLaN2CbYwRZKArdNyoVRZLgNTWBUO//QDi8J3tkT9FVBe2
i36Q0ovn7sPa4kTGI8/hkKymwzJolvhet0OskKQ7SUuuKUEe+J+GwVinSIa5zWVwYIR4Oxjho2ul
chnQlbtxewEYTPLokqID7m3eUMXYEyz8P5hJwlGHcaJ6G2vGXOWz7uN4dsP729PUKCw/23HFNO78
3QIpYemajVjonFzKcGhFw2ELrJNpbrB6g11B3FRHq01LvG4JFm/eWIVD54dIMOYHyWPc0S5ICh3Q
G+tKf/DSVUE7AqKuYPhTTdbEenniIvkl5lI5w2zXknfOFwTDgAn2grodQs8fmL1orGrqy/1w7SZe
2uhvDTouwUPsw2/lvS/Vo7FZNg+ghVMgxh3kKc4Nx3mK2U+hOiQVWNaHC9tCD2zH/5L5WbO8AXcJ
cGFkUEq9BGsoHv1yTZbiFdc1XrPP2ixiIkrqoa58KAhBtQ2vONg+5BlOALrD+xivw/bFWZ3PAEfs
3UZpRt8E7gni1XP44DnOFIyE1Wnt8bhOaOuou472z4WN/61z/41REDFpN/4m9/IokcQI5Yu+zuNA
x1uZtkRd1BDm8RWV/e5jlKS6KbM/JhA1EcWsJHv8atJDcNVbrGt8SFNZqA2ByoiIzL6w5FPbL5rt
mpHTI1LUpc3x2lU0j5HEPEPxpmxB+9qMsmfI+6Cxo5fiIQsqS1IDv2W0WNfxii3B+5v8jpjDzUpt
/sVZQYoP+zzve6oSSc7okcz6ChHLc8Um68hTz+L4hXPHMp//grNpzbYZNGw9INBWFHn/9DIM6QaQ
Toaj1riAYevhpe0sDa5pJSStjBLnZXIDFjbH43KF2FsC8skH1sq4chjOxBhN9pvrnQPjGw8zsHFd
1APHc1FWBbC1xEefO6F+wC5Csd08DulOQMmwu6vTS1of+8gLWaIChfyFAajeISFkiVxTEx//7svP
xL0hKvURqbPQNFlhyuFJMJIbIcaY9jZCu2ByUJoqpHTWbUTAG+StbIZaQOyGlbmV7zVQgm+Mh9Dy
LwPyhBAXAtS6581huXEXj4R7PNdotdKytbcRnBNy4BkD4cWAR5eWLffx5+f0u9z6RA3ojL6Zg/E5
LMYWrZZspwAls6TOHHs7qMjZlpcdglNqqI7O2LeMYlulvGxwgpeI6AqNCcrXH9TblMRl8npjo6pC
5FaP9mb0XSvBd/bsazu1JeFgbS8+We4+xuhWNwyJrZvmRceT6602SHFKQa7o+4PtSUIsFAoyFlDU
O8OLiDWVu/MGhjex+uPBl4I1G1zim86ezYsGhdYXdJpJGAMT+79aZry1Rvx2Fj8iudYeN8NQaEdp
Z/pSdL4AiUiNQ73mtG15Vh6x+H1ak3h1deT7habH+6GDAyvH2w/ReuDEH3ZQZIKrBFEhCGdz+1/X
HAlTJbarW5DXG81i4REY2Sb9OeevEdrvqKxns3LO27ZTFLQQFM5PaS9rlz76DmdxqYSVa4xHO1T3
Q+9S0+ABO50xnRCozg1ttHPhamSTiT10cKr9yHM8dm5Y2JgAH0upe1wpBtRKrSlsKRWw2vqYmqIX
i8JmwXnQkXeCvsxMoYFTSm/tzrs4MoMNeAHmwIM1zwLQ0OWxfbMoJn1mieKP/rFmVVdBj27KOOtA
BosFVJTK8HfV8zCjWVWMvqdZo8yXUq/vBbBnvtUMpIxLfhc3zaEfA14Q006ZTfeDcyM/gwTjNJPi
YSz2QPxp4T/pWj2FHZfBlQOkaou9h7GlbeZTJjE8+2moeQPgHKgOqt2Kw+nf9Bozvd11845Pn4Ua
nphzlE/XHMZBnEIqJf6gHaLZJbF8NAtit70M2qE4iIhnjPrluyRCwiaCh1nAs1h90+Ep6/FgjvpI
aP9Ckf9FDAD9zqEMf6WEh/gaTtxUWuxKA1aOn3RVIQv0AtvxwrUtKl4DK7yiGNbkdIiO3E25ODB1
bzZ56QXNiVqwwl++cNM7natjAtXP3yHMRjyDvX9DCI0A3jneOwIQ3bNYcNP3AKkHBNs8/jyLO5zl
MIgerXHtY6qu/mpVq1oGq4dnxiv/Mc3IKEaKoA1p3nqa4gnHbdAvModae+gh6yZTN73yfTbeM1a3
91plBIBmJmgUE/G1sie/+NSEOVP2wnrNB2SMzHW61aT+nUBGy8SEHB2R5NOP2Bm2YCksaXIUxQWb
xzJ6KpELfgwo1PxPEm7f8X0db2bf8/MmANV3DOzYdYCWyNB3FHc/lFD7sabnd6bgXjEJRPYPwfrH
UEQ//YrEK35JM2tK+zGMSkXnPTSxuHKxJZ2cBR/HGQ+dXEGBy42xAsh1Wp/mNT+0qPuBsteC/8LS
As3YXYWLzakEKVJE9fEJ7vkiDdUEoraco1wHp/BQYqGEseYo5AmAXtQWOtHgRDyK6tegTU6Vre+J
GN/RE/tI4a0Uxvog8Vekinh84ZHywPvg+fhrd8XO4AYUAr4XZjcOJ65nAq/E8/ECcXV4kdSB8t/V
ww8iBtqlDGBsnpE8YbLG/pGMfR+GygJw5McBacdfhw8/ylUO3MK2BRAJEL7/y9GxTkyMQCLX3L4g
93Ky0bE0wOOgP8ww89H7P55jTqRBuSCHeaEKcofyUZJnpngnC5mcBld3NmdIgkaogbC5UFW8RqTV
XQWbIWDsBfkY9PXHk4H/QFp5j+WTrQXHIc8Ii2zxBnLo+X3CYuhbbyY4js1CBBqYfMQMI/XsuW4p
lJ+NNWiwyH21JgCunSO0Z6AF9cgOPr+zsubEwK8Hm5m5+an8ZVtB0yVbmMX8Hix6wPfiaXwWOFMJ
Fw03vHQcg1elfKUK3vv0Lq4G5usvHJIwYZbLFkE9Wuuu+7XiRRcoiRjskNeifMof8QHGgqSaXqHn
cVvW1BD9QQ39S7SDdYevwMGvfUuOLunrIu4KyuXvLj+sgPlhW8R+uzwWjLhTXBwxgjppyTHGq06I
7Um6KlcsrNswWiGe98Uhk9NaIOQ7c3Ks4TQcvWe34/WydvU2rocBguP2tDn/+QaUpIXjvXBLPiEw
IEX6sEfRWhXbc1y9FvlUJ7N8SLJ8cOtje22BrnJ9OEEeqvxi6Y6XDKQtN22evp6XQvoiCykNdMxI
U62GQqDUOr/+qbxRUPk+7gHF2jV1T82q86THpa5P0DetLYk7yWgLDXv6/hZyO4uot8vyNKMVAdeS
vjU61cNAG/PcdTnRzjQa+biQtxHTrDC1Xxr5sYBiSt0+FVlFPfhJQj3Mdf+ji8HE+9tvSmiiq5nB
AxlN+ZPa6H2Ud06Kh8JtsRR1D6aSurhV8M0r0NKIGUWFk9AmieFIRWPj3OOa7Ts0kEyWzyu6ZJUd
sZ0GLB5OIQy7DDxadzxFF+vi29RrOSN3N0nTIQAiCTs1oPcxYt+6OgoXpozeyVMRIr/BlJZZIUJv
4DPmEMRZczDV3aFGF150jcyIi8IqZKcVOY6YBMaazL8tXhtr23671+xBfN+lutei81LRGOAYRIRG
pNIuKop6tfAvGb4nxtWZm3YS7BcDs8PiuYlEUnVtyzadjN2KKeUfJOfkB2zqB3KtTGxkKflyaW4j
EBaAvD3ywvaPqtkoOu+yq6eu7ISIiXSTT6DF3yVT6JdC8Ld46kcaJVqVNWgZ1XPg6jBEcEhyGuTE
eOmceZRxi/Cap+oXLcSylUdqC/amiFLaJx1FJ4UHj1XkgAVvllMq3pVmSa7akwKnIE35+hWUJ+TL
OJ0LHOIQGDsTK4PfWjH2G0+3QpMeYehSNQgqHC7wXbEJdDudbvjC5D2R+RitNUtaY1ZmGcBQKPeN
jDIBu6Mbh0YPyQLrHke50VoK0ZFHxevVq/IpXbeL35LHiHK2e7//6Y4DD1JS1NUzprnU1MrvUxXn
/1Z9KEuO4wzsh6XfxacdccGNG3IWAy9PGtUhxBEEQlW57GRGX/Fkbu4Mp8D0cbtS6C79QeBIwipq
8FeRGkUjIN9Fbt2KAa/hOmlYaiyWWQ/zwI6OsWAS1n3jwJ/2S6BdTNMp7JkUunZuTvSbuusDpbjA
FG67If6GwOLsrAZTX/R+iU/I37yOb9yol7ehKTEG+jGq7vgdr6wHCHfNDcVDQNHIiyKxaHfjRt3W
9801VGmSFQNN/Ch4omtixsDE1pwZp4FKk9p63zYCQAF61mbyV/VUeaU3R2SJUHPxfE/AF+2bg/zy
EJTRhZ2lBeJINnd4Yf8fo4TEZ8qZcf1kZkgTN7lII4qIB054F1gUYrkAJcO8xyF5WRRTzHvHMLHt
a1AKet1fkwtI6SSdIvDD5iSi7usZL4PYdQPMB5x4PcNwE7rm1g2O+dguCk6k6S/6Eah2mUVQx1u3
+pVIE/cl/Cnnfhl9TdeuK8fic8dRKUYt5RM0bcn+0Tsf40TuhX99WmXXJtQwNzwl8AXDac6e4daR
jA4bWtxOgcT9BH2bUlGOoS8/z8TcKpuCrsnoWucO41xXFeOlbAn1LrT5ARrQVi5DknigtDKh7yY4
BDdeXKGu3M25lokwjg6VFfV5kFF/xmdKG6YuomrroCmpYYr4zmP1VwFK086plyE83PLP4RApfG4d
cXj8e0v4Lumfyujnn1VRZXgrZ3QKci4AJvsen3SykEPrsQUHYVyOmibBnh48t8ymbwi/u18JlthG
/trYoxn9f98r9znB4P/pCjwaJX3yt6dygRBH6s5gWJT3nzP2fSUXZj9/kjXGyqLQ5cJkf1+13pzk
RWF3t9N1rjZymqrAfU2LMp4nyzrT5nhGcSVdnNUJ7AYrpo3q1nDOndDXGBbe+IkR7t0C/hXiPe9l
7ep7lbK7xMRKF++7irWNt+sKOg9c4wPJ+JwzX5z7clmVfwKSjhqiFrAci7lQtRb+1PJp2Vu1B383
H0M91XHZa2wfec/jnSPz4ypL3H5yxAzhClEQLfij6gf9/UtXTkC6OZ7CvEHeGJfzxu9l/NouvhFb
duU/4ahEcnBc0WFOZqVbNWsnLRI0rkDTO/hyKj7MgAYngvmRPFp8UCrOqPNJGb0ToQNJwULmewLz
Wy24ry+7KfLVIGcNQibMjOY7hH5++hL5xRPCHm2260eQ2JCTWQcF2l2EyoCysdhfKpo92gmAVhIz
0iOed4Rk+GwXP1zIwH6S+TVKyn7QULMBL6YJlnN/mmVKik9oRaj4AOtaKgfADRHtqVPUJq409kUt
f1LFhxscBnkb5Wgk4CJYmO7Q/u5QJWIqxUv+AiXmktLIKgdH/WAv9kY6Xdw65pjAsoGjZvkDBnN9
4gofJBfwQ1+SeJSPt0SuJ7Pz2FJoI1a2dVVsbJVbDPgwuflTU21Yqt6ZNZ8+tbVjg7+O2oVn1452
M2xihOjfAjnse5Ek5W9xv7iFaUnp5rQRx13S3EsTETaAiBuwUo7jxjHV8KYqjsxddUqjqg4vAhet
X3JAi2/gY0qdApxjYBDa29hin4pRJPyUIIP4wh7t9MDJOEzSurOlDTIUT+g89AwOozA2o46TD1T9
wYyOFlO6VRfReT/qQX2H4VJuxqr2KWg1bZSy8j2prK4X2IaO8D1b9FFwuV7m501XugsMMbGco0T1
J4cUc+OXVgSXeEAtNo+V/LxIghQYURLSFYtxZy2DT20arlNA5kXB7d2ZUOoCtfoRjVMIWgfZqBgS
IS34r+qIhzXBdUX0Qf2FWXILNy0yH3KXgah8SqScGvyWJ/v0fpZK6YcSIo8ZllrOhBjkMWEpXMma
biqR/2zhLhRcY0PottPgnG9iLgMfX/YOUuG1mVCMNS1iccLWsNN9kRm6MGVa6PFqPavgPADgX2Mm
dVnMVj8lxajiUtxv1xDuRsSS+0mXWM4YaLEA7KU7I1aveg+dGUIAhHrV+xOY8gIg2tqPoT3b7mBG
pV+7hFpFcUcS/mVbsLz513sdwydpJeLzF5rqTL0Fe6bMQc9pmcrGAfMNgTuG/whHeHmZCSd3hwLs
5BYHB+Uhqic9mTasGg4IMXoxaDQHrA1kTGvDARAJCTL8ZYeiDdb1rOf562LbLLnOuIGu9DWItSWF
aXxr6PTzvtkfijR97Jvi0vEKPyKBq5uADQQmz+itEazaX60Wr/WFBrdQ9n8LWh7PnVfusZN+kgNG
a612BnTuGPP+5djIc++uvOr0WTQCavN9taoXtA3KeiOjIAtrhejdDt04arMY7Er2NM3lNFbEFXGq
a1mLbEOtWob2uuPglgNER2gHw4OJ33iO2GvKddW4JzzPDA3E+EHnYPOEF9flArV+Es+RRXgRegCH
A2fbJiGm76WbdtIkFMtlfGy43jYdMOctxL3Pv+71sd0efzYOgI8GEK7FnwcD3b7Fgj8gl6UMOMIU
++9yjMy64hhrASBqCd+17gRqYghZIBUu61NuYhIfpvMyuBcOkdZvTy0wow9XhqkiWVuwUpBKFWrW
2G1SCpSEHEzqbyJIdjxgp9+TwE/VimPgPx94/iRE6wKvYdlYMdRneRcmoSxDOc476iMfRkzX57kg
b8/N4buModYrH/QKQoD6Wdm4JXTztXKPbQ0WM36IXXPrP4dX1R8aCchf7uyyl53YDwzKiakEoeyE
bKNHUywwIHCItfO6fpzIHhCgFLkozXyg/IG8MyWuwST6/T08vUY9I+kdYI6rIYbtmTvbgW6Z/LSj
b6YisuYZodByb0GC2z1LkPY4gU6VL8COKcy7E+5Suj2eS5GngbNu8rU8uH5lQzvfwGezpIzGmfir
TvML0Y2F2/nY9s3QU8NG4Gt9OVSBwDl3cpJzFU+hlLEPzZPZPQY39S79UUJYN88LptJU9KjMhltc
+AtLFQAc5IfvEz5/1QimRKyP84rht7QH7Y/OLBm2utadhMhB0unSzBCjwJy1QXpWV9bUIR7Io0jl
MNIkSJ7FvZq/67WQOHWxuRIo7gUoGyS6e8LTUJqh/o+QtLV12vnWunQnrJ5d7ovMSllrETRUMIiB
nYrL3MfBpRz+mKJe05fbRs0CnRN5fCK+xKxG1DnghIh9QMAJYbqO5pvN4sUm6grKOJXenVOJjM8h
2xwAW+n4pLe2vL23hcexwwyg742dSDr6sv12bnaeud1E359uDHLTGxg5OualGGhCnqFllePwHFY/
AWmTpiCqHGYOqirAs0isccTiJ3AhObve2YIu9ADKfs1+7P+QzxRc+OKgelKup4Yw/uresCLhtssw
8fZU8UGC0h05iMmcthi0v7K2/tl0hgcetfg/Z7PSWbVsE+cOuG7/8dJzKsdSBNgVvP1hu8CE/j+p
uBFFLVgCPRYw4vJ8sH8oD6BJSGsSBPNV0oO1biPbg10L8khMc5QMBIrS2kfCWn6MJ0L/XNTdfdbH
+Xb5XOjWIM5RN3E51Khj/zuwa3E3O4s7XDoUO3xDJbwei5ueqAxpfijLBOW4A1WJlHiTV9Oh/vjn
aN3+8ItDdkY4o3MnZkz0YJVEoGpl8IQjm+zZLB/9F8tT06zWYGyPztLJcsr/Cgaxdl/801BLNRIn
eQ4oTKkesRnNuftmEgEd5wntC3JZMcqoa63IXwcJ++7otDKbX9xEUe0xmvs2o0e5nCO3U7lluPG3
hbwaQ5AaoAlKzBkKMtcWUX0Fk4XvXcm5QFOF76SejKT9kEfKCeQ+n2iIBf30PMH/rfYCTLkGXIgG
bakBPBQelLedko3GCTGMxK3DoRWXC89jcJVByzS6sw+cKqgdEFR57ErOndonwBpKMMP4/j22fCcY
1QAsioXr5R3YIhsmlhMfNFzrMrRxUHPzd6EsEVbyxsStwT3dME1MBDXlP/hJXv8P7nTWHCNDNvzp
555PLztv+BDuajE9hYbkxb8LoRbbZSconEpS/FGl9QguwcAALxFJGrRW3SZWRujz1ICDnKGnhrZM
u9C4wV3mCv2zpy1Skv/ZfEHwNkJHU4XodwS4YYVoRfMT81hstW8GuBjXCpWRYROVV1JV9Pmxb3pK
eoAFQI1taBfa03hWjsNUFP3/32ndwTTWfJlJU8xf3m/LVYvnRAs38w5e3ho4CqTT+hfb87aPTDfO
zvHBOpmGbVjPT31lLNXpwHVsJbqaMqxjrL5wr/93v0B4DzhZMgvWxGcKnzJvVqB9NLCuLR7Fjmoj
PQRDNOkfUPaLDbmg113TzfYgbaxXuOF5oh2X3HcItj3d85IikSNLgusN8wBN8UbvzQLNBgrZQGBz
SUka2JsfuEmEQgHC9uRk7aYlhSSWk/1BdL8UnEuF1tSJwJEpBFO7wPRfDf+yXsHncdcTq9Vrs8p7
6Twrwrq+clQIK9vAenK3d1bFQAXqta7uHRwCTzDMZAeHgb19HrpZmKg6z3zCiwWkhfxlDncw2xhg
VNV+L2vjZJaZsYghN4fpeH0g93G1eCB4A/GW0Z+pyO6lUWQV7Klwa2gZ3/EtuH3puhPRtLS+SUjM
K9rrg03+UbqEiJBxiBuonJCDKLgn53+X9f926Uk2QKym/qnPtC/JjolWVtSAKsmR/sT3NlEo7v1P
Z0ezIieRFs9oqRhvre586B8qTmu2oYSNX2o/jI/AFQYBgRshg2DoJYqgxORTKezqeRmnAyJs3rvG
7WeOz64MYHgDfNkgTrOv2P6QEK38UcuuAvCXPAR1chgtk2rcDL9scfwtp5GGnhynObY47/KwPfSN
fNTr9+2xblJTQ/NmmRzZ+b484XdB/x/VjS3L5HyN2GW56Wuk3XSaB2bcCKacZZQbrtTFWn1SOynr
uaVnqj7CPRf0DyDx26zQ6JPRPXa4gOFpW+cvDmJlK8Cx2V+YDGdxYDDQ3NktgQ1/P3+Ta6+9uN0+
uIyXZFNIcRH2pkHQMYE20VkIrG24Uxb6ZlGf7fVBGmZDznOTLLr7E5UHXfiumkb7Tuswq4bmv2wW
DnFAz/qGLkgdlNZjtM51wjSPNfc8CRmMuwr+ollGRMjqvWLwuEnXg22jzAMtdCneOm+PZoQjGnqi
YGH+4ZwFo9OZRff2Ai96LdVoW39RTWEB+sO5YJjXDqEwJ/cK+44R2lr3pFzLfEvBzbhIN7YMpY0W
bAAiX1YB+X8wFKloU05gvnM4dWTMXLiq4MRap4srjtc8vEzmJIvt+FIwhQSvLDkeKU7yHwd245il
6aPOlNI+f5nKNaqCBnViMfW0zwX8vjck0TLeSOc5QB3sGATxuZopETWL/KwVxJVcopzSGNlt8RSO
ErNCauKTrnxXwj+vfB9ThymJjpe1greC/Xkxb1FyAWM7Dl4J7kFqhRNBWWJ+hI4XM05CXK/4wm7R
XdM8+Ob5h1vLmorKehH+RK3hvQZAivhXSF0EmxQ2F/wdxr9ov8LgxqUMrZxxS4l54Ge20jK/5yDH
hz3vz1VBQ3xlv562kjUXrfdRUwG5ZsGq6deAO1qfJtClfC1E04gAeY32Y+Eqvv08I/mOLt7AEvr1
YsMMaciHGbNMPszw1IpFWef0ywmCIlCctvC83AxisWFyPFgv/gNHFjQO8OoM8KAypMmutZGHFmlN
4BLbEdeWl+jcUi+KoKDuCr9unCWVeZ1iyyKqNr5KVnbjjl3JutpCzZ02pRKA+zn8RuvR1tbyA7pZ
4Nl0DDkR6w+bOEnQXZaP+o/x+b+UaDhMDqiRhqjaJLXWNmKpn5JEa5dt56fGP7uc39LglV4biqOu
/QG2DrQucVr3CPwgIT5NPbnNuYcL8g5KZMmzPidsLw1KtorxpldRkxcof1PkxZJb1RuQktM8EoEH
fiupUj3nZ42cAfRzDfgIQJP6QaCjyiUO0++1ZuOhweyp01wVRvIpiDUgwL8mvOZtgHOoSUg622Dt
tOaRlOZWVpd38papTLrYY8exn1cLhw5Db6+kWGUjvAhuKCGbg01QRqYB/9GxH7VzWjE0QDkaeDLj
jkLAn4QBCp/V11DzNHeTUGcWMxc+jU9yecGnjM9spLuW2U+MaDe9SqOOX+EmZI4hZa6/U4V/qUqD
XVRWYSt/DI7ci9QdEjed2hid0Q0X3p9YNVCYp6j7HasnZ5WflsXhnPRa5JCxjLWjy/525o8BKUo3
8bbAi4MxTBfdHtEWNXOmXxpwNby/8GlRXMaJxUq8b/HurVAWEjNWQJCWMaKolKGtsAUcpMMpVgkb
cCMEvOxsCZxNH4QpsLCWF9F/wWTeaWwovNvfRcwEY7uZRtURbq7u2DF5UpUmWs9dyaAXhARBOicg
e0ojUyhsZsxDKKRnaD3MSjDBatxeOcrPz/b2XYFn6O0bAok/NBKeK3Biz/rH3LM914lgNUYsZdVh
I8im55PoubWZV1zuG61BX/gjPEAu5DJxDWzvR9Ds6F4TCCoD79ASCdqH994EYOQz8NYRQEC3AQJ9
0aqtgUNIygDjyCYR9wQKKHf34rSq6lsthkdfBM/aYd9uK2kWhYRirmuVBwNz6qa/MRfaOaLEGcdn
2Hnn1rppfnxMY9Kcb0kQIWYliUgoclyPEr/7Uomt+ykvujvwOVD3rUECt7hbm2OgXvm2GSG31e4S
FX2vzfNOWrMyMd8FKaHjPkLIm/WGj+W+4OaIZNMrmm1uSiUIdBJQrJOihX+lKWFuWRQRqfny7uPK
jIW017YKmdWdWY19u6vJFFsgrXQYL8Hj3TgQ84Sp8b+k6ICN8MPU5oRT0RbS0lLm9WHee4do2zAa
rsPp5yQ3my1bHc/0Omo9e+ds6iWXPLdSCU2OOgJRhwATuT6UVwJ3cMVmxjVST5sevB7ij8JWDLY2
kY17FpvO+8uinATEGm/9NASQMhsG9J0qS5lBLKuSO7SRxH2LbJE7mBQGbP/FL1j6Jb/2/leJc+Ls
K25PCqveLOdLSDaoeAvBfVUnhe22e9ztHho6iXAPY0retbDT4klOGXRCFNGpFFOnLIGKEaQxJqPU
yxkyEnSMqYityO9pMhoXtfVysn9om9ziZlCt3TNNV870p4MxKXKWcV9P/jm50KdTWuRB9TwqCD4v
83d5iwSovcs5b9jLlin2HWHc1oQ6SVF5sFf33c072IWbL0vNlbemWzeX7U5xaxFtHIbIsnBOrCrC
EnzQlkLxHIAP0jAC9fcyeQgkmmdoVOfJsSBQZxRv7J0XDodVFF6qTzmTqZ67viMIVjo/Jb9Ycghn
mzivIPV0SGjiHToAiM63kR2V+QNmTKyCnZJ3mjLo4S1A4VL/LmDpILRSmOzmqO6cvtQQDEpdQWyB
23gCnbIzS7nxVvULE+morvfyv7DW1O8OkezKMKLemOMwIsPO2iptwBPl3wh9gZ1SKiF8fhmv5bBa
Y1R8eejqzhW8XaTDBjDfnUBE13nWqfWpQQm7YN1tlfWHdqSVQG9Daiq2NbTiCzFJcXtc4DlL2aPJ
fXdWSOnOYrZQ7SH8TaAkoEGXySsE9nrgZy8oLI2APUFziz5eEmmKUNXcQO9BborR8bSIYOELIpAp
R0UfFAZycu3YF6KLNMvG2rjcbNs2YOPv47siz9wcEvub30Aobar7ZDarZDoXMGqW1VCUcuVONgOW
rZY5VJnjqs/WMwfs5syjHmT3a1c7ho65Btt4plEBG8ygJe8isfHEawfSL3rUgD3Ncsg/G2I32UkB
Iv24jxPxUp1ER+Y/gGgkteDTyy5F46g29qqc7UkJ69gv6beb2Rbwy+FIqV05hWQwFMeKR6o8SRp+
PMbORlEowcp+FvT62A9Cql0N1P2D4RI6VEpdj0rI5yR6F16KgiekBa8hGi1Cu3U9S0v5bW49YLxi
8g7IowGwIwpYKGZq2DkoadGHqkf8obEwqlMIqd2t8hUJHyNTaaSVY/x5IcbM4crw8AiyeOX3vm7n
tr63QevoLvO/AQjudLPq3FnWdNachU4ipeDAkZ8VKdi5orzkfq+jSxc8n89mm6P79UG1+Mr55zJs
CsYX1wLIf1ztacafoda2cZKQDOLBKsCQSBq2P3lNldXdIdk1h37F267ZaILsXHXZ245na9cj5e99
V2eYqcuE9u1ufctv8DgK0/VlKSscFJTh/yGku0PSQn8xbeu7zSU7CL1jegJscK0JCmFclrZx0hdO
cfZ7HOQ3AQwil4/3qMoVG6Tf9c3diUVoQzEJuGikvbS+7H+B9MiH1AEzG0aWedIbGs9SVktaoJXN
IT7Kp/3Wi9Q2QP2Lda2Uazd/qaW8v5nfxogG6prnuecxYTHfGUSJVizScVuxLXKO7AJEXni1fV1Z
udQv/Rqpz6CeiZSrGBfgfAuxSqeV4iJA0EnbnuxnwOKEQcpbHO9lNhk8OGGKcWm+uiVFtGV3x/UK
Sxr/BsGk5akeIlKOoS36Ww0fTFG655R4y4dKAZtn5pgOD/HLlNwB4MMCZJhgJXFSL4qnMY3tfxZ7
CliwP4GWTRf2Zq9ZY45fXPUYjlBvGHKvEIIYzOFdwKJZy7YoASyW9iKGv0Fw5C0HxpnJJhSpWD0q
24tizPS8so3jZczjlb1okGHhB71ZJQekl6SmX5HgLQlL9CsX57wSMopfqZj7+CB5DhRXb3dkb3B+
Noa8fCQWnENmMJHxSpOB9K4vHHhs6sJpUuifZGqF4cbiMw/J9t26gWP3lP1IJ76C7Snv/HLbNWPE
blCxkPXb/M9OCu9mg8Y6ASJignvPQmRx4a4kzIdXcVE+FG4JVdyWGXPZ6RFhoHhd1c9l1t0WBuDa
pAx4PwqXZlLTDO9Afq4+hnQm8tPgcFkmMg5sn5uKc9Ob8fAvjjOw6Ul5KstlWchwXNqqfEt8Jckq
csmnuPNkCXd0qIwlMQsVzD/qSW5VuOb9Qa2IQ3ghn8lJ0L9ovKOUQoA+K65pQw3Nd180ZSBaYuWI
UDXFDJ1LpBo9PrlXcQNB0SYPMH9YwLiHwjl0h9mvV0o26ujF5KI9h+CSnnsyXqUsOiY/BeMYe6h4
GT/2Ge0TkKhLDmN3zN+A9oI02Zp6NuSpB6LKkF0LnGahRxo9v0179J65yX2lIaLseDXFVvuIbt2X
0PkGzkvnkLVs3UjMtcdPNDSLaLxrF0MIsZ4swOzl3WTG/W4uVYmZwIwC21dEjD6TOE0aZRLxVRog
1TlmKrIia1aKUShcfP3iOwpCiuKpg5dMyfE+0EZ9XSNcHTfj0XlQEc9zKyWFJqn120/Rl217Rrxi
NJqWjWShlIZY5JpGlkGAq8mQaUCRxPa+P7i4j+ubrmYisEsVDv96JROlaJqwcFqcvUzvf+Gumhrj
U8WmSz8MzDoIaXCUa8b1vUt3xoPdrUztr+M5TWQxmuOK5lmGpiZqL0+EC46NlbhOldgnZa3BUXgs
CzqRD8zT1piEYKV/IKdKosoBqA7jnpcWVApEqpzATQiGPBFrk1cfs/ZKSMphdenVqxE0jTzzGUOA
WQafwBkLrCLaXgCPnydB1hE0UZO6hoWwizinRN630OshHcLU+s3OIDyGveKWszkF6YcYu6xq2Vbf
K0GbyG0ux038Y8ouPuL3lLtA5ZpbwQoGrbu6+1OHzvOZfBnnpXi4nxDSnDYaZ79VlMn6JOgzjk3Q
D8M4zraPyEg8Bsdq18IP5ZU8l8Mq3rGzeZFzGsSKqsYvyG+nzn+Gc0BrP7I0Y5Cj6/u8wsvJmzSN
F1EcDGRB7sBXD1rvl4ncxsbRHJZ4NroEQwAqo9JVrzXCHm67hBDJV3ebREzg/9O83HbfZPyvhJF/
q411raThyB6vAHxC70OGbWTdOWAC8fe//eoL4/1H+cae+b8R1TCxzLLzV38HoBeJazmtSKeLrNtq
dK4ZOJIGwGvh5hga+/35MCnaz20ephiRs1cL3QusxEIQ7wWzQ5lmwMnmbuLH4ZbcenBnPSGdd49Q
/lcXLIm3JLjZSEsWof06kHbKLRQ09SJAJifiQmIICHmVXryAIRhgprD1CziDf5zjlRich6FQo33b
q7CmdwZOVsqjOxUC1L1nwGrAHmiBSMJnQk/otmzgYnoJoJ7jMDk+2STOTaHuozPtET8fn7g6f3K2
FNuhhIXEn8ZGMxFexBG9ZLsPeJIyNIC9hgaJy5SGkl5hnLxRTLb4QO79cGpH3FBUJYxtqMfmhw/M
fW7LjYUhGYyqKCveWzCT1BfEX4ZFkNVhbzoByKeL4U0XCVPyj0/rOYceESKALfSe19ACfkpU1Q+y
uAHYdcWHLxII+wgmTDDRbf8SxjBzBgeW5PZpRv5dTlfkeWiEsbQP9jlS2g9HeiEFg26dlrb+M2M7
AxoVJ7cCH5iVtxXsqRgeLyKeWzpt3GxT7nGkV6JpCh88lxttDDV0QKa/6tiFnanP5+KKtgaCpIJ6
MzNB+m/z29yPWM24SguIPLndeT/mUi4qXE8VbMClSDHs1BXlB2yLre0Q4zfwMZpNzBXHUp1U8iZJ
5s/E7G0TDOJ5EuRazNWGm7958v5A5T1w8NM9JyNdmq7DtSrsIHdk8xtQur51G3P4bqSGoZ+yhDec
UR1Q7HYiDJefwu1Bccg/qo0be82LD48KrWd0feHARGEtoaOeZCpV36sj2fAHWbEB5NrPNmGg6Z3Q
AwNHBwkf0P/Qm2IZWNgbWCI7otIlt0SAAUaYE1yGm5R1yM5338MTrR/1X1y7VpccGndRt5BK4KqI
DZWFxQ3zn4kOeqDjOKijWP/PbJ2CfgeXsQf5Xu8J3Giea5kQX1F/ZKCR4jPb1tHYE0hWM12WeZy1
qU1Df9a8AlW7GlT814TdLr2PwyIrMyzpkuWaKr07z6eUVH0ZdJ7G7G8UWj/swOBH0jNGIDF8JyA/
tqJBeG5IrmejjnTLOfuselVEFgvHMKaG9NI90RvujbMwjp8ksrLFl5PBEtRRy8EMCoONCtAp9EQw
EUMDfa5yVy+zBKwH8PhLAcuvjS8diorzs7iaSfUltwLm9Fl0dxDBlqWG4Ge5tQGouTUx7VgJlmOU
CEYB3T0WtPkxjquJe2a9BY685DD1K8KoAoBzluvbXHLsurU5bRURu7lK56JSQzX/+XUF6fageLYE
C4G3sWtILxoIDY5l+W6zS+j0jndyOtQVtBbyP5rKpkS1IxRrBpf+WATL6bt+JohbP00aRCGYCLwa
4LyAPNF5dl+wcM5UwPiDlkfTryv4vTW3/Q+72oLdT34V5/e4CozwaayXhONznR4/M5oi3L+1xc5a
ztdRaxiKhCea9otAmJ7fA+4AuBG8oLoA1eiKupR808aGvbcpa1P2v6Vwa4/OOHD8cprniPkxqRdD
C1vA+rQ3U42cRmjlg61/pWIufn0OvmDrK7rCt8QzVXUXt2kdc/tn81wd5ax3nMIZ5gqTMFQli8ew
6ufarkYKOAdZQmhqoduBJj6Bu9Vwcl6CugRHUYY14nR8qOQSE9RqHfaJyZnPMvcQ4r5W16DLakl2
12UJK+SeuZ7OOExOqpXhmW1FC12azqaPUlxim3vjhGAsH28Ckoz6L5lg/9ZFyXHrezOu6MXxPdUO
MASAi9UbrInUUx1XysVZ1b6uwYlpdPt1mkBRDNVZb94c2FVRCAUwXf4OrFDZ0EvDipIVf74zRB/9
2LJW3BU8w1MOYQPEA2+ivl33UB8c639kMflzgnYpu8Yw0QtjJHgA6K/Va6VBpogPQiSE0i87DnMy
BYl+CZ9Q8fimAfm0Q5RIC9IjPgbMOrn6K+pREQ+TYDSKjleHL30LMQZICTaEbV/VD/D+UjdhqNuE
LyvgFduwCY0Ln4wKIKLKDz9DM21jbvAR9lr8Vm13S2v/jeM3jRZ6N0mtY9Inu0agqy2QnvBbwEgS
ewl1Z8MA0X53p+LmBatgzoMa6xnTi3jqjWjbTlTLtPqtUmYmFvldl4CrsyTthpsxirM3DEMTKxGw
vYIrm8ggBhM1WY8mv9jx4fMsIyb7ACM+gWgHRfrqPQAc+RR8g2uv/PWxrVgQDZYxQptzEstSvZbE
JM9V84nDR8ZcIJ7nbxkG37cSC0RxOBBTKm93e8/pfWqKoYrs3BUMPyJybdnLBR+0vQGh6eCyT6FJ
eN+dHvKqcSb3/LhGDuP3VGCwzH3jwd1Uc2ULFrHRFVirQqURy/p69fsU2rWSPhu0D3Q4F+hhhAZ1
NEIA5wsjc02GXPjuAVfvAyJbThUyeKyXs2jmejM27Ch+ymlz1v0+sOPXeAqnr2YmbeVF9mrHogPN
MK/GtaaRTTtz9lY6mS4lHC0SIUAPIA3ltmQLyBp6qLWWz8HLdYk6twZH0P0Nb1N8Q+PaKIyUty+N
A2FyVZysqXEqPczhTcVdRG79ltv2i48pbWVVOPsonD061RT7qgCHBKcLPR0drqgIhUzpxoE8tY1y
O1euZDRjYQMlTYg9uvBWnHjUiBBkhNlPACGRUeTYlxzmPqrHjadknhk9Dobz4KGjTr1l3WAHEgit
T0c+BtC5X7HlObs7+J0syd2NGa+7qe7RbgOwGDqAtNwWF7QTzjtpsP5Kgt6vs2tPMcZvPtyJxM8C
Vq+FygYpLsvBSY9JjZ8nrCc2AhJswhh9O0RrvDe0b0WcU9nbEbcKD6W+WB+W2mqKxKSL+vADtSAu
ULvA0+NpknQn7tHVdpYE7WGolPq6Deu4j4VquKpgg0kBUnfJ4uKzt578asd5pjgNDN/fNz9PSq8B
VFcDD+gr7nsiAE4t9MYBZoRzxTi/cMJQjfHs8wS9xGt+0UalAHSoHZVIyqXMFcRj+WVINbiLaPgI
pe/FzujJ6gmqdR2Ld+9G6LbLHkD0OGHfbHkfI6IPrsD5Jxiqa77KfXy0F9j5vYPEmEKsb9QLWSCl
Ki8o0wE0xCRHNj6tecEb+KzIqPNIJbjyMY4V9CHx0yvKrxJp+aXomKPpoH5a2M+n+Wqm+RUCHA6e
aBjLtTp6WwRBFMC/3kJQm7xSLZXmcx9sqsvOxZMczbfJoH9rXJytUv9rqd8FW0+qJHVmQiMfBMHZ
7rvHpT+xQC9esu9ZGDLsoOjNcdLgsksISEi6LoqMUQN6j6/d7GUzQy+G7ektG4jEsFiKX7PHsTAL
UR7T7cRn5TlqvfUcpVFJlKCUIxYaI9QA7VcjJe3XdQ+5SXP4BdOMlRSEZSbqsWI2/hnXxlSDPkVa
JwkcChD4xbl3Ti7mc4ceQIc3UvniVw2ihOHeN3I+/+2yxV+rLVoQBA7J4QnBCpCSGkNGAhbfj3Va
knaXwKH83dx2H2e/MS7B/MtRKDE6MYRcL2yDkOWdM/DymYZ5SCBabnCU+zykFTsnDBRA7KzLISuw
TF0CrboMaucMjtwJpdeHObePhJJY2QjOHm9hFYaICczCfE1gqgkAo926MA5SsQxS62j9coqkCVh+
C4OYmnRoDMVJtvh/JgoXFphwRU4O1b9cU8j0ZlSm9U1QgRdq8rda/aNe7Bqs8ppopmB37IwmKEJ4
JCKK180B8vD2Wm6r+j3TVkda6PwSEV4UFSmVekv7QttywjZgH1Dueh8wpS9sSx2ehSIatzsmi1rp
vjJ8YAzdCf653odFasHHUFNQXSd+LhaAGcKR5n8xUBnvuxzyrLTc/yjkrZ7wmKUwvsXDUa5K3wHJ
D7PuDrIZRHqgoIaRj4Vg+9HTRjUMWaNT63s0sU1OkXVaw4TD/ibebXrIUvY3u9H2opq+UhAohOSa
5drXKPUqyLzNJZN94rx9IHmKYLENcQPlM3RWzUbGrfT/qL8V1M6v7iSrmuGAc0WKvmUqQK83snMz
sR/bCYU+TXmYFfusqxZzbrlQFVPcxmp4XRdwoaYoljcIDnDM0giN+tSoi9nJQF9hNkyCdi9iWZMd
zIdDwYlSKdZVms/84QJJfYhS+dO0qITF+PaxjQPjRIBsA7dA9CSpDWUHRKU78XNru9Fi/JzEbv2h
tnuGC2HPQYH5jyLwH2M3TZ2eOMV2yJtLu/Z/kKk4ndHOJWleJzH6gOhxAMHs8vdjFZ+XIyeM6JUl
vvAMfLQ16wN2oUze9wx7BMeR7zyX8A2k9oED3pu83578+vyIJStei9qWrkjoB+LBjtgEpfX+mqVl
CefVDrGWW1S4qhBivvol77NZWWSwfuTi/OsGea7uBReG1gS0DfTPomd4DjiPxQwDtnnkDiooNLEr
BWhGImSoVORxLWHt6blmz8S7gPLjd49cbF+yjarlNjg3NJse7Y8ZimXkG4AHWZYje3SMiHXRnGCG
3Nzdddu/IJielF/aexnFl+Tir8nGfK9h/COERAkJ3fGAgDSvpf1auvT3zR9YvzvClwH6BMmFHQHz
9/ymLPkDTjx7kz5NTNntVCfn7xDuoRuqA+sT3Y8ydkjWe7uU52bQk/wtarAegARaApYZv15rNb6T
+l0TZcN7eQfUEeKjFolAlkW7ExCcc8wxPge7EhzcAP+UOsUMBpcOgU+vX+BUV1zyirnvzvNbNRVX
3muoZvA1UYeg2C3BQd+d0z/joyojwcSaKxzD9IuC5S+l+1cePebNFU6USPyghCcORFKw7sw097kL
pcGZLkcGJDlpwh4KCAnXqPA95uJGslhTFxefVFfauWAgZOf6DZhuBSQsvaV3Ld1vemBUYYBLr8mz
hswgyRJ/fLUvfH1l6Kzptq7WCHyAvk+1fsbpig2hiSBLFveR2kiD3lp6IIMfKj64OwGWB2ucHvmu
OQ2VclzHHpauBATjsD337NDm6UnI79IXW8iGBz1pSkTK+1XPUEL6LdwQAOhzQnCMLr91t2xSvo7Q
4fJ3FGLDiuznE/B4dzGPbTA5s7/eqw6Nh9C8sK2yetU/EHwj5d5hfRlIbO94BzsOSNbLD/Ot6Yfy
FjowZ60PAUZsXgz7t+Zc5p+eo5C0LWJBcWpS201TamgvFO9UT3SNESik1G9xAjFu4FgzDLxBjZhP
DUBiwSwpl7PnjPXuOKqDL2Yh6ZnzTc/QKJcFYFQhZSiTZiiQQ+stQLy/AnldEDmZRYe9fX5PexN0
e4XVPEtFB9g7KtPiYfWqSVz90r4oe6ukydjNB3+sSwgN+fHOtnzVozvZ5hjLVJdsYg5wn5Hg3Bd3
wjNMJ/U2rkHvHfWfg7920RRW2nOG+cjZgb/big9v9e0JLA/QGLm0XdG5Opml/qzss3e5ktLewVHS
Uzv7vfeO12KL5bBLzNk1JA3PFIWC7du0lrF8c/TwiPXi4V5qIKibYvswSifP3qP1J4sB3ib6ayqU
P2QKuXASg49xy5G0x4tq4G84yf6n9eocqr4YExcmRYIoVPrJ0V5/jUNwR3IUKy1N3SUIPyQDf+3T
7cxkZo2cQBVkaRBTj7SpE7opwnMrJrvEP/H/akEV69dluMn5JWXkv1ZBaf6TVmNC7+XofBISonJG
QbtgQuseThHpR17OwrZYk2x/Lep0beKlKtfnmH2kDj7E+mAeZBeTEjo4xGajGdmr4GKIZ5+gnDYL
js6sWE1CWs4v6JyLcnU8ZKd+8YjA8gCEArnLMS3bRGNA7a5NyJsM0bY8E7KEkZSHbeuCO3h7gOP7
bohDkoeBZ0MVFneqcx4LCwR/4QCfRUaucyWVxSc6OAextohmXJi+NpxdV9tjxSgwVxE9Tq6/IFjU
7ZNfsUYyX+5oFmCpZGuKsgcb7gs2WUfl1dgUrcP8Nb8xsbUqmHY+wEWNY7EI8SShy8Gx/pZiHGFk
UkbHanRagfiSL5H0+J7XP12PUAFUmDYlq6Y3HxxX8DDoBQBZcG7tZJQ4F5WHKcv29ypabZ5mHlvl
sWcOgHi1W/A1mIXlKArLUM/R5qzR0Taf46aw1vMH9vuqgrlQfbLy+zQHqWwP3Xmakh0Y6vNIfQ25
J7LkwiS3+RLr6UgAkVHn8WjuKw7QR0lazSjwbJhd60WaVXkjhA0fSdU5Pb1gj0qA5Of/s/8nylLo
7t3PCwEh/fERPS61WiC1pnU9sFVZpvOqXAoTxtQhRq9owoOnfzKvHssqsbTqysVhg8pC1VihzyTE
BIkz0DiUtzibw+9eMtrs35dbmC2GtL2zZNNHFx1U38wQwX8LgZ9nutTYng2YjAqU5L5X3bEzGk07
atAGioz3RAr3jMewrNE4EeeqLJXpZ3z7Om1GCzKL858MnFCq8wEBfqR/vGV6lUTx6KbaNB7edtpu
Nn76s4LWgfVZDBNevqFxMvgofEyWDIGZxkZ+ROyLJaAcp9VISkGPFAUx/GrLxFpaZXOYtr5eko1Y
IyEdJBMyCNbxqoYJ1tVCTKCtJkXyGEMlkq682ZjmAuUY8SXXMYZsQ+6k4dMGX2NnhKxqBcc8aCPN
UBahohCJo/3uBlGKbf0pSfayoZ9F5qziF7Bhj6n/wsY4szRhPocAMs4+G+zpoFQ1hZ8Yq8E2ARnm
3PLW8GwGIckc6pKyAdXh+VpX+TY7veBKC7cci6B0Woq7Dj68xRlALP5CQHQib9nnknlyUIstR2H3
au7NhHQ7ZS+P7+KVo6Ng4yWWhzApaoMTQxIDVBXRlbsLr/GPxUhmeJ2GNzSulADgB1TBgUW1XvgW
sswJyH2Qw5PcPAUbcRNi/HWNzq9v0k8/MqzW/MjkNKt1XTEFpsopHhLBMdTksqGBO1zwIHkyqoAC
fKDOY73AtB/VZViTKVKCirKUwM5PRydDEsOV5TJjN0kaIF/6sNF4j7bQh2uP0ucpIoeaVXqdpprb
eaTYIu1SBA/7UgoaA3qGn93wlhuuBCHen2jN23e+9AmsYL0veAHTjusSrUhoj2jfz09E36xz+kms
vpRPghKm8wR7kq3Dy0F2lc3Golaxm8qZUR4odGLUHQXvpE4itA4x608NpVehiY0VFnNykt8wlPiI
H4znTqY1l0Xnj0xsGwxwCLNcrCn/D7f/Jau7mTpROcS9tVQ6Fp1CQnBtSjW0eaDCxfzLXB+GBGMO
trRmJsGaVIh5ydoMtjvH8QlUskUi7z/j0Knm/6TUWMZh3cVrLdjLPeRxnPFKbbnK9mqXxp5MZKrp
C00cp8PLPHKmwEGAf6BiCeIQK53ZE5uh+ysBH/bkiA38JFd7gFNvWrt9hHTVP2xFh2Gcd4u0vKIv
1t63BL7D2a7pibzMREIPW7QFlpYy9tEcIg2FpHAQ9AGHk5/Oxv+7D0tpu4TqJk1eCwy8iUhUDSXy
UABpCN9syj5M3SlumCQCKPMPn1C8vPFi4noUqB4XHRCjchY5iS9YdT2e3UnBkTHR6eXdLywVTcv/
wYLs5O8zk40PzoioIw7N8u9pm2n4hi7vrZOfq6cMdA4AyqtSA8Bphy11rBMZauQvjPreFfp+7RT1
Cw93gWIfrv5mRwDO3zwBV4UixdH4IkwV3UDdmcYKQaHEuZtGZpxC/nbs/M3+m0/Kbmyy8gVQ5h3G
Sz4+lo4lD6UNnrKnMJrLaugWK8kdPKAoSKbYy9mo9c/rTaRRNtiAbvhLBya50sLRIl0Td3LfxupT
aAYXGbTNbtiyrEvNb8ahHvyYRo7BHtiP1UCOEY+LzS3ZghGRpbtecGQGj0P8Tn5RJVVOgBzX9LEu
/KHs4x6ClwqSHVDbXkmfMurTSDjBe2DtXBjJ9RNGz3Bh+YaspTGKJSaiprkdBK/yX9wH7CBNI8BH
gdvO8FZYqMegTjhz1/Y+Sq7A6dAchJYiHPgkMuCZ53MYqZtsyqPMOll26MKl7SwPeYMjn7/r5MAU
cRP4yJMbzRk5ASWfMs+JozILuJTkPPFZ6JygNB54xKgnp6GZAj7kHRrcwwsSbPOaDmh6bOctBiEl
uDdaA4uMkReFnrMXNCxDPtrAuLJ7fxyNEXhUyN9wKRX4yXagIHcThXEcUOLNGcSLlEpHp/USYjfS
p/PeBz346lfnQkXd2jDWbAzuOTtn+8yeZdJc9y3N8f9d2yIIe6oaeRZi5X9spqo7fGcv3OV+D6Yu
k0v8yvu7om2970SEVIQoB/g7fgesgfIBwmRd9K2LVtUEmYnzk+BgFC+azVbS7yQHBVTS9lkptYWw
NOKwVwOpVaQ4uLx4XwcaOFyYQGyAvDWwlsRqc77OPBBhj1rpapin2trelGDXwMN6Xm9CLQ2Gx/gj
cj64fiwT3cBsEJgHCPXsIivGJMWaed9/1R0izHxd2GOSSigeUJyadrSP51ADZDr0yV625FKS0Yzg
YbiWkVIC19dA5ws665FNwln56R4XgbRmQo9Sn9BdB9voN/oFcP0PO0eM8Zh9aeK1DQh2R6uFJAl9
M9OQFPCGmIJqmApGfo1REZ1kcO1luh9NXnVU5Hs9/Beuu5fCIgGFG/MyNDHmU6ed4AYap8Y4kZms
iWAl/GDGNgiVN9y60urTYLuf31dHvWrta9vxNSHUFScuCXDaGQoH7u7k5OFo2rba+aqWuymzhW8w
WfmgbpOLWrHVEXtp1UTV8+dk5ZONiG4zsNWZbROpMAWfy2+8vTUJF4UqfgGGV3byqenQfjgEBA7g
7GedX7g8Jh2HZSa/cyzV4Bn+vA32fAvGp+6r76+Xt+W+wtroRIOyj19Z5fmHwTJfr52G8FaWskb1
90xvERkgDPe9DJDtcvIxgtcTMnxVinrkrrmtmjaYpVyflTsfl2mNxeAqVqca8gAsw7zDfCZBGJJG
8YeBt4pWWiZ9OXlVzRiMdEmgiWZSzKkPVsju9xZqBARJ+Ht0lUCfEWuFKve/VNYid34RIBUH/Vb7
L9ACoPi2JvG7wXTbzDp6YVVBtSK6wygfotC6fRtqVMiy9DZrJ8mCH/eP4znX0Iz419Tj7/wtRxnn
0XPXGtVsodYDnhbb/UlmAsGhzs0CdHHyKVLKixxpioaq82St27+eka7350ddRYabZUaQ0/wZDiu5
KiHPGyN176C7CSzAURT9PiSeXkyKU+lHB52NxbthgexW6wq3KM/0iRrO/YM6IF5O9GqqNWZzm+Lq
qq0I9XHqPyB1dQwv2ZPdDYOKS7PN7RDH+IOh2MkHt63Bs1JSZIvmX29ewGYNTpxwWjdlAP/byFgT
muPTlnXnbL6oj9joVjv/xCwJV6j7Dq5OHiFV4djF7yqrc7/fSHrQdUy/oTyt72RsItl5mC+rz1ux
jQoJoK63Ijpd9JENVBv+SWNddEgEdzK7kH2NiIvztv4Qi4DD0KN1ncsNiDcjOcGgawGiaCdpRLno
v7wmla9H9+FS9up9MOpuLiXqGvXqpZmSZ+mJucixBTV1GXCYPgiJso+86Kf5v9eVatiCmKLa7/hi
5Dc/pAI7KjKFxdFLA7XR7yWvDlhtChv55MLudYpgxNXCAWU+EAw0uzoPSZzPAmPKQ1pZI+wgRWY5
rHn6yoNrV+tCszZMQlR/7criA2LbtlQNtajclhGHCAZO6IaZTd9q7JR7k4ZGOLGFJ98vRWVE76Q2
V5jXqoc9em57/uQ4VKyzRYbkkbP08gF1qTSalSfEhAyak3IaBT6J7SmzXqvNYtEbq+xTZgTFVTmC
dc7WC9l6cRrX7fEdpXtANkf/AGiRBBv3ZfMTs6LBAmk7Jd3ww+R8KARRRuH23GH7dH0Bj03YUu84
qIg8xbl4IoHLyum9DiROITrD4engvz/GIB5BCAPsbNBP30jbRUzpM81uAcVuN1ybqXb4lpLCHSJ0
NEugRuQ+o6YvyHm0+feeBmLyR9xwzWVTtT+Eyp2ONRxfXsDYUmn59MpgM7eYvWklYd2IA8CnJ7N0
PH8A9iN1tEXigy9FMbVseAK7kwH8xNxxycIdvQVTea48MoAFiNWXLi05v6r8HjMGWkHEpakF48OE
KWvrluHNQW9oyNtlBDPbtHY7JinPDVSaXWrBaifDDP09vdu+RP+/2jsJgjhcZWdsY3sYPc5KRag4
+Hd28B4+1cQGOVK9ulCwkwAX1wnCtxe16jLqN56ndMh/kejPdeBc4J0umEF2T473fkw7F8rvP8w+
X6z1vUtyN2iTkqQmFRkJYSlRywxBIIgPbLZphequchXHUeM3KPagl5Gov5BSAIMC3wxiiFd/LnEi
Ut5hIfA5kHgInlA/1PKRb8gjfG+J3/PcgOu5+0rpD8Gr+UVEUM7WBap9Ls3zeK0It7kNqBRJMMeO
DtbWRcSJk6+EEdut3RJ7CSnp2phj3Sft9y1+DZdrwZjJKzjJ8mXlJ9IFMVNwhcL1XTAopnq/gUAf
aEgqc5hzOVHrRq4VOhQzExW/mDCbgehQ9mRpZb0pkDHjyirUj9giyye96DjS8nJmg2U9ws+ETdV+
FunNQwmEj4uMp4Im8dPHGw4QePuEYULJriCJD2pQqG5QLE2a7NRhbrVr4YEAR4nj/edX4ygjWmBr
mICp02VJ+Bq7V5RjqWhuRsEu8gAwttehrEHxRolPJLU4eNt+d0dQ2tqIeyoHr8+MwEurN2RewCjJ
7wa7rfjzYhDCSEaoHZTS5opg7uhw38W23ylcnyFg8zbYRHxHsvQW7Op4YNjHgA8xXCkhjBee89uw
xNG1/cFKGSRzMCtJwGmhLhrXRbpl4dilTqFZf8aZ1hTMNkreGmGyg2FuRXSLbg8dY80M8WfsBgLO
moh2e6385h2K25KI4PuQ6eQS1rQW16Oqw5VfpaO6El0Kg6AMl5yryzEy8bVj3hrSeqrH9WizwvRD
re6B94Glv1j0CpiBqcM5XFIw47YB1GmIXeXrfdtFlRJkgXMUClkHCYgscPPJgDFbo3vaet7ZSEBz
mLcqsOw7tyE0IGb2AZ8Jb+dNEWYJirwo4odHvnrgYWead83b5IvVduy/Ozn2Y3eW+CfOU5dsAZ4N
EdASGEfDfplWvmwMsfTGQai/3eGODXXmPHdzR0Wdmg72RZ9Cc1tRMRQr1kixdsli89GWv2b1N/Sd
MnSRK1EdYHaJlFsloJIIoOC9FFNuG+oDn8D4aETc4EvkLJwmZYN1kZ2EWQVLesQ4Cd38M6bdvxGk
Z216GRVEn5WAQn/NeaXEr0vfMYlAg9ddlLY0HRVbOczHtH6rtke6sYE4qc1xEhCo0EBX3u/dGBwh
28VP8ysPB6b7gfr13aw/P/2sQx8LlyRUnlmMhSvQ/YqNat4IbAB+fJBSv4VMO8zWbRUoK26qA07a
v3vHgYvIlG/lunsy1D3EolnWZ8Ya9yYmbt/IyF6JaJl7H04UdlXVqZSb/nZ6YgCGwYvvhqHxIbS5
9G3xS//oupqepLd2T9EMcUYLP3dHTaeqY6a6cKIyZolsHQRaiPa+NsJp0czlO7bdwWrycfiRucbb
Y+UNhppbTJ9Zj0xVacxlgGSpdCP7ExAUT7gz45IZWeD8AfiQSwRNo6VYBpXuINk2BanwBNFGCct7
/RMXj3YYb5DR6UApZOGypiBBmxJg357Sqxq156dBV1UwRQ6VnmohQ1nyD99IRjomi/S66LgDhlCX
8ODpzz2DK19UmYMfZYxJUP6fFE4X5fhR5hBN0C6t6YxLtOm2uun4OCD7EXCQwLz9ViYvOespRCPM
D9GFIvNRI2wFOYGnq6TYVlWIJ3ZqhlS/jhijWB2XlkmOAllTa9JOyu+PfIz3lftHj8LGBasJ3OSg
tYixTk2YZ1oOODo08WERuu8BzTMerGRGCPPLlk6Ob9UH7UErK665PLWO01OydP2ARqM/We71qOci
7kki6Tcce7kiHbF7F1o4GU4OiPLp3jche2M3t0M5VE0A3457ZmQuSdgimPor9oPvIHFFokdkxrw6
EkgZeObAA6K9CEpZ6GgbmBNIaqaRfMrRS/5dSNDoq0OPQRE5s/2T5Zx+DlOusYLjWLod0Gguass4
mIGBcPI9BtdO3BNCU0w73VLAy98UI0YYI36rDKUxFnE5ydTu8XUbJ+wmHsadubcyhLLxcNt9dNWB
CbMbhtceBZQ3iYEgojoQk8OlUCFZBokbFBVboyL0ZXPeJty80/c5YG+QOoDEWGvHl/4TfLXmUxB5
3rIky1bNuXbv8QaV+/W1wVnZ3eVQ8+6LYpWOa6vMwP46cBi615lJhcLdbhA6mkxor1F1dLKpVG2M
5ujoEdCPHcjZtKbyH3yCL4k8kdTkHAISPti27oi8ap1Zmzd8/39fVqLAOSh7MJDN6F/xSHJOmgVz
CV9yvkeYD/kcbIYN0IF+okjm0cZmUnFXtghDbHhL7WOA9TUNEOU3NsI6gS450YfgfE++PPlObFNl
Qgec6Uc6Gz0zP4xgEZpAfoxhC7GCb5H7sRALFFUDWkgoEmq1q2puwIzjr66TCNNfQm2+huH/2YIS
/PA6V2ucpW5CNxLjSiOuH5GMHNnctfCwm6xBaVlKApxezROaT6g1pq6sOVXejxAgjYuQoWpX74od
8SNvma3SEK0NFOlL+J1nxjQZlepY9IYRZl6MfBKxdEOQ/rYlNbDevp8sT93v7I20SxSiIx2FJao6
6wrJTJq6Qbk8cKZZPjWGf52IbJQv3r7ju1mAdzDvzZms3Loa4uGihQ7WmIxjo70kRsgs/37mxMDz
xn87r2JKvLwaLs+o/q84O3U9cajTVJzUZEMtkTLGhCkTZjYQfBzO0XTWURqHWbkt34Hbr7MxNaVF
Gd4pXq4BoqqnbqzUBRyvf9i7NvmMinIEEliyhLcAstZF9KMUnME8iHI9ZUsDVQK5HvN0EbLiNG7B
Dd14q5peUJGUYFYks57dRA9xAIhW+9UNnupYpUs9osM7IcOynOT+Uhd1Zxmr1Ki1O7hApoXIyv5/
mgm2HKpuhjARuejDmzf+f7swBJN3WxbZK3pzPd6OqEUHnxun0zX/+AFOCEG5eGSEURd1DW5vdsbn
hz2TPR10qzucxT8JR3fb/dJ3+iG2KL+GA1SGrNvns30vs9U9ylx9CazyVayqLO+eo2xV3cn0bl6T
KfiG56Y6qO/Ca1uWpu18ue6GG56BROvaPD9gHGiXFCcSkghvLJZcFBL+X1UoS0w24sDazD+Ejd/M
9+14aJgirxfyMkxY8C4dM5nWXTwPDDjgj4jYNAzeo/tU9nfsDb38GQu2Cy2VIab31XPoW0jnUdr7
O+P3ItlCsmodB+TLHxqN0n8TFS6e/tb/b3yrN0dJ3gBuUAJ2KLMansucGcAIegNUUJXJ1sORuvUH
GmfH5koKW3uSRS9ZBDFGJHSQn+bRyCI5qrgZOoMrgQeFlFlNKzbHcdym/RKI6FNYVkEGFQTF4xyt
Hqxr1QL+nypJzeQ6p6qKTC0QMFrmseWfqYnXloYlJEKybpNkw84Py2S5uFREvi8VMdi0foq/395t
P3aJPaR2fuQnbM/1ThkrgoqMD2TDxl+CFCTq7MqsqdL+u3PU9xV48Ecg+5MIhCE+DMIz9+jT+Lzo
JIV6H9sxcIHzFqg2I3xkox163Xk06cals9T8kvtA11bVlRT++k2NlbbdxAQatjbOl0TK98WzvgSq
vFtsrH8QHZz0o+GCfFy2AQqkn0NCrQCwAUegxQNTDagmS9mrJwdDysmRA3KVSjq1N/pm1Aehj1hY
JI2zWcgPjsRF12upQM0fVdOYLnPSCbCYNlNDyoniYnDc8yJ0l4nHcLnXFfx+xuAihI2JDsbGKWHv
ehMaNUauBh0if+S43/kxrDE3uTUYS/MrGng+dyINNEO5Po53nIrm524PuaM42DF+t3KC5d3c8DBi
K0RdY22us3IcpY/Ydqa3kxKcGWerxTCw6PeeaDWC5wWZ7YoOD92BnSIkxu8bMuPI5UvinQBPhJpM
2T+mwSPeLmdVBotv+ivcDqkTwKNUvf0GAXXha/p4uGfyx4aYYPgsGi62uGOiiM3xpnnbs2JvPu1d
PbPU+C4Q/J3oOEbJ2w/9OYWfCnMi8CKiSDl/4t5h6GyCc+1aO67RifJJYsBslz7wrJCMu7+7x4Dq
VcsdeUfiXkmlkGkMPLH9REpTWM8VuS4SdV0C/yd8AH6tQY1u2bG+x5nmz0WaTXLDKdrpNmztidoh
o2efGNGb/gm0h7iMiNkjEftCDE8LKyBvoowD2qMSjmBgVX8lVT5p9ep97Eryc2LbCI9yRvngThA8
YA10hjFMniDsYT4mx+7rT7i/ruvgsYj7iW5Vl6pQRmgGoeWRffSW1b6hVVaDlSxJ2hElvtSgD+h7
5AXfzRJ74zbelSMeDrvaxDY6v/jA2j9jCHYVJEI/drYJuXNmYANZzZiw/rUOuexKbUjSoPig1OlY
haav6DIpDfXOpGKHBC594DPrDJUaesdhTC3IXDLWx+1pNV9H+o5hC+FyAPG6XwB53HOHr6knl9oK
52ju7/u7+RUpk5JdwatIwexoBn5v09+5s9ThssP+/yBACucWzi5A9qjDAm3cWzCDytEOtBTwR6xk
pKkJsrxz2ldSC3j9zevhrNgXsqxabEyCZvt5f/0oCx9s9KZxVq3OZ5fBI4Lt+QhqLVOzT7MuOhM0
YEeE/nUvCNVFQE99uh/EoS1C7czrQ8nzwD5fTUvzAr6GkWYIRvX0OnEL4rMxcY0WEq9lUSt7GXVH
QX4KaPovNbLokQQGTGfCBcjhtKwYj55IkCJizXZqh9vdilg1xidVlrOYoYgL17Hd0shtL/Dhqxuz
0eEN6hH9BVa1ho5F7Qw9yQACi/+N2qS6t5XtJxJMH9UrBzBHc/1v4ynzFhN+Bkz9wqsX1hy08lF1
7kIiyQoVZFqSqKcDWMAfol0EYCOD/JlzLPCIdxlCSnH8TX2AIf1zxKcz1jHZvYzY76I4obU+gXRh
cj4rhhQ9ZPVlkxmEXSWG6FZW/KajUtfqiWBos288oC4m22N0rTKmofYBCeMn8nGNbNcZwxmtHvHm
JmHdFw94yBz1qhBkd+g8Byao+MJjPeDn9H8biw+PcnC8rc0bneocf/L5mkkMMpUelFzw5dWRJzNz
IYhw9sPFiDcLZ0G5LaWDF965sUwpQrqxStC2Lj2WKH4u2CPejNZSXdX47ZzLBt4uhVvj75kCZihK
PQyJpdnEzp/ukVsA9zsz4FxuSlaCZylotsUxuM8XRQkQauPS7baYwwFV9ubu77Olz54frILc7cB8
ZmJbbCUBb0ft51KKVH6wpZO1pSUisJGr/G3qTdGKwpgSI/AbS8CPTAxrEdrX8a149t+UgHsKMCs3
KevRCkrOGcUlNQg5sa5lLphtFCiS8hcUwMvC39LtFLDd6tG9xzqKI56Te9ByMGmeBGXucNTGEwq/
r2+x/TAtNqDPLN/sSsPuyUP49mD72qCqR/SQrXQzNGqbIHnvgs47T3hnh9U2fjCTxbCu7G7Sdl5o
ad5r4+SvsaOBZxbxAYahK4n1z9PBYB5Npq/4kNvoqQz+jnb4ID5+kgM9Oh7NlRY7ECQVN2woRynM
1zIdwQQgXT2hu7SpWMmNwlYIBRQgJro6aBM3xqiXTLEW4d6FAfnzorheR+a9oV33gFt4iv75iDAE
P/RBY03Hpgzv4/rLw2iE05EoyFpim1DSDfH+b46/uZsf/F8o0lPYExlgEYyBxWeipJD5vg4nEJHk
7R0r2BNpJq2YS9pyjoqo/Zh+wmnk8D4bLMoNl9aA5a2dVODq5PGCQe8GVTtuasMR3ioRBfDo7rNd
ODvza5dEIAe2RKdySoEPnU+eBLifAxLnwqvpYuyWII+ADy0KpkUcUvrhtGk83EBcfUdHOn9lyKCu
Y/HRSGS0SDqsc+CjL0LSQSQRUWzqNP7VGXkHO7wU3Ps+bddyKR6ky4VBkmoiwq7d9O0khpnXf1Yp
3YSMtlNcWd1RPuTfArM7v2GyNihSXtab136MZGHm5C7lnep/MZUMEexcAgOpLSSpmQPIJTBtB8VX
DYtfU5xub+KGlnpV/9zyC+RwFw0tJvHNOUduQY7TsPSS3h/fdA9rOnFZFoakAdpsspPy4mtUP2hx
Q1QRN96TJsE+Gw8FRlCVN26wHAx8Oa4rerbFX5Of+NnuEvfDdbdLD1ropvTLeEvCdQM9DQsQKzt7
n3QP1rwDAPNaikBe27cdpNGVyYqkMXuBJdA1tnk8MBlkkogmQkEm/b+XSiEY4vwZ9IszYIj8j5tI
0K7Qf6Ci/GTYlH2hQoagRPy9z5OwAePjxsqPXTDx1Zj2XH+NTp81FAOEGGfYqAZZ1ySBXxvfQAtJ
6AimZqIMhztzkHK9ZGYeNwrZVSLq9MqVuvNHZtmJP0fn+KTJnCJVtsNBNH3AxZsW31hXvghU5W3L
9XnAJOplqNyUtsmlgjN0mErmZs3SjpCyqojhE0haSWZci2mvLidkvoxXkoh4D03npmIewE+qx6D+
wRJMuM5YZ0htkhe6QOWqUJcQO4naayr37NcVgQnh3ApRu1+x4wlApvbUAaHnQu0sRp39i7Zo+0vB
RXi49CdpxPhYM8bEKDV/h7lkPa2dDl/0qLd6/aU3QKZQ5bPu4tSWoulW0+yDOwo+BxgMYvAL7dAp
dpG0XMty1fR3uuaeIoEb8R4mhaFdsVaF+qUTEYIoVupXPFJ5oiWxS6Oj3SA3u+LuJ+yRFAb9k8Ip
SdqJfOs038efxqCfHt3m/1bI6i0Nqf+LyjhDQ8nOGrdweWbXzDRtnw7zo+kHbzUp+rxXRYNqDHzB
Qh5pbd+uh6RXo9KK1NS7n2n/fQnyXVxFRpxZ9tWNuFtpMAKjryPM5H1E5EtccWia31I4G2u8T5oe
p2Xw53uIjIgYiE8oMzzpfYEP8zw+JdBpmCYhj1Na5wfNBHLzR9wUWg5npJUrHwxJ1xcteS9x7iEU
MiYEO3Pbjq2pJAFUEF1ez2nwBXrqqHxAKmycq+sV4hEx5e26VrCCsXXYihTU8lOcQkEDWLl17NtG
tzQt2zsCCYdow61HgEZXrxSiBX8nt8065y748xofbf9M/zDZCdk8f4cODQch+vpz1iYLm1+KvHHB
goT2xUZG2mqmtAOtu14GifEecmHkOhhMZJbroPbbBTKabrE3gmZ4vLI7xOj3oIvZcb5YDrfhqVWY
HnQz2dLxBki4XzepeOoH68iciNlUsW5HcWdXKaWbK8Iln+DH83nrvkxT1zDv0QKYMNMrdhRG4rga
MJp8OO7/ZYIF+p1bs2PZwvkJLxj6ngZORw1R07eC+sTdFHa6PZSM+5e4b+G9jNc9oF2M2bK5Bapv
9uBfC7bIxTHAedvbIIupFzJ7TaKSJ3ZbhG0YgRL+MNoDEKw7ZzPYd7gZRuTHTor9u0Id8M1IFBsf
XUeH/cSIwdbKugJgTcf7e7RKEPsQ2luz5v1YJYCe+9l2aGFsHmckqWLbGf/YH6LZegicoDcuBWO1
M6i8YQ/HPfDcDoaF+QUdueu+2Wr4r6CB3b3oXJQxkX7AURDZ/CS+N3ywto7eVCtTvGDZcVQLh5RZ
Kbnl1povUQbAxL6xmrLVPsSueiJzchiU0sWFsgkuicT9JJcrQfP9mCBDJlfxWoy1KyoqbKMlGKbH
70XMNpToxZSdsZYSAtRECQ816VIUWSsNu9vVom2uJLlotWmlbeF3lPQ8Zu4ISCnAtUwp8g297h0e
RIuf/Oe18mPQHTUMgyKvfMpZHmB/fymI3VH9Q491KNjiGChoYfcNqoJonuuMy4XCCAkd/qKKhCUU
7yU5T3/Mqb9oyDuVoPZX9hO/zu2op4IMp3N8rBTa5vA2LF5wKzrY08NIfO3LFwy873P7D8OueB9C
zoqhsu/7+V0Ft04JRu14N0gqUxmi2ilXpAwhGOY5ii7T2zWC7UnGvfn/ih7MWkDGHAWq3yYPOMZM
7IquFwQYkXsG53IsCImEM/x1h9A0J1txBRrrF9DVFV9H8cZiKsoA7CLDNROwpU/f18bXQJKZiksI
kWXA9uz/tswk8dDYTl/W2bUpwzu12VoSdrK++bub/QtFoZpnbp9EZgxBk0IhTTKnl1lupkr+k7NO
I51XnGpMfgv5d3ew/gw0Rcabg89DIXWaW1ze/LWas5FcUG5AdOOPe5opE7sdfLdhggDiOV/y8XlM
qcSDwGBDH8nwDzsnoc+lPkVp0xMFbmePTE638WSP+I1wjNW6v3gAvRrMw/r7lza4yi4jS6N7+oLz
oa4+RlWSecJFNzdmIz30nEbskSrXaQhc5XGMNvhWfJ7XoN5hdU9wk9xHPlnD2w6rgrTHOZyfFKZD
HIpfnDp4nY/XbBA001Tnp0uUN1tLxYRl5k4L9/SNYg9OBk9Cas3XOU1QW99+B2LxSrvIV7beUqIU
oIsmYbRBO/9Qkv1M6Uh84S8gmA0RjGrfhU8Le59bX/t8QcGo4nVh8kH7XF9agKxxAJi93eHV+LZR
BbkgnqnVBrJYVxini7wRpqcJnshf6Jxh89JjYFyY1wuFvGYU0Z2/FZcUT9eO59jtKlJgpSX5u0PB
cWBC1iEYJiE8PCDDZjk/Y3jpHBc0IN6GKn/RNCgsVBbOAM5Dko9lH8SnciN/UUGvlgGtjji+J/Hu
h0CBjrJARWj3hZur3DgDOqA+JEpvzGaqHTaJTC1zkgmQlTrp6WAUfqdapuvuS2fRhrDNNZQ7eJD9
hHyvK6sSuLdkasn5P86rXPVOrSnOZKDjTvNZRkj67hLYBmjDOQpTIzfTTlAuDAP8o2AuUu9/upQr
XNfI2EFtnfal2XnLszMtXeyKNp8t6KNLy5hNdwhtHc/v9b13YylQAlJPbBH4rcmiR9442CPRDOdJ
TqI4AsQUYdMq6iro4u3b2FXGdH0Yv7n+NrpxhNSYIoPbchJ7KXms8ZTsuTs3b5B4MGEZyI9GuIDU
6eoYZKn25zJ2ZS6R5QSVxPLivCHq2pjQo8zoy3ICWUfDazILpMMalCcXb5K7yWtSI82YDqQGt2VQ
AIGrH04zTPmbM0ekQfzyIVH3wdQJPtoyvmxA4jhVE2KadBfCGO+bOdr3CsnBh5FouohChCpOPsju
7N3ECbAJhIty4oU6R1vPpRSQ+GtFxiKYlwEHZmM1PIu/NG1BEq+KK/IhbR3VnVc36wVptc8vZ0DW
sFr+kJOaWPm21CxKn1oU0cjB0LKTppm7v2RRdnd3hhH5BBFL+W6Br7/HZ8k6lJAtk75rHt6NwkND
YAjCarOiaPGy62HZFHLVCBy7ge7nSUFqmyW5z2Wkrl92onReeLEBs/zxwa1IIj7nqcipkcrxYH8d
1iKUU8wJm2pnYllAvDw+uGejaRg/l4NtdZIJwJpt9huo+5OmthvV4CX9Hqss16U6KbipMPNUZFot
owNI0JlB4vzajloziEQRGJ9ypmzIvc/AOddkKCZRuI2OIXihzk4t2z1DHrwqTtQtNTS5NfINqlE2
K042zzIW1oVfSUV9W10sokdAXdmUgCwZ9JEy3BLjcd6VhLa+qBfLxpkRFkqRiezbqtkXWUm0GHbQ
1gsml73bf93rnqUhe0fy8WNwuYwbxT0ILBBlUL8OAQy45dx3umhDuGLU31YWCgUjMfJ332ayje/3
Sa3eLcnA6r0mycc+9RM3PxYRIve/CNHmvsP0YCVSrDj8ZghnLfLdX+wm56dYiLSwEhoG1UU1spad
bkAeTccjX62FTK+8aumsQAzL5aSdngJgKes/JCAW8pn2wacaxpl1kh5DXF9yE4ibIur9y4LcHCfI
JcctpSfgxS7Hot7OMttJd2cclksRVt3/Jj2liM7r4/3adlAacXGYgT6FORp0pHd46uRm9I5yA6kh
Di1cEL2n3UsCiIe+14JInUxL7DWUK7vyGhINvvB92xwBavtF/EEFs6ukRQxlc9e+PfaARcAWLwP2
Q55At7FOmkYUO955r6Aw6Bk3V4jyEyJP4FDBgzJnegeegmgoNwriqn9+Z4+R5pdI+9uDnBF0nt8s
InAhNd9bv71O+UI5wfBaxMvLiVweRHptF8gJQcwBmKrHj/E+vp34kD7wExzzRcdhiDvGtZXavC0u
50FHoCVl93pYSjWO2dQ6ETBUV/D1SaXKTWvMydFbTd+LXXRRYjvsQhVGzs36bL0aN3J7qx/R7Nre
pBytsaLjvWq4xL+cpC2WUD3XbGR8k5q+Lsgg8tSMCoF+0t+TcNEmd9saI0/rfO5mhSiRKLdx8VzV
3pn2HSaDzNljKsmm3IdKlF3C06iPfeyMCRf+n1jP77lG0KDGpmRnpJk9MRlJ70eLkgZVPaoZaIF3
wzqE036BAufdTevrO5fzzRyEN7jI+NFlHKYAg8i3jiBPiy1HDW/miGA5GdDBIDfpWalcWD5TnO8U
O21W7Cc3vguM+mXAUaHWJkqlacosWpypxzxIG2EESMLlG2cx9KzvxpuFQxWt5WOiAHPLyW4mCQlB
N3XuD1WK/anOGH8yK29SgYSICUg2cimwVZcUvGjnF51zaBMwoi0UQsQSM10CdDc3X3gBP1DXmHpw
nx6hPAEQSCCFkQSfjI/E10Q5kQ2hxtmYBSGfSUU8g+T2nau0SnSVG69ic42/tVSunYk2821tl1if
/aIeO1zNR7HstukmSt29WmOPsQlQ9fHqMgfP8HMNiSJwaWWBKHTdflAYg1TP4MsZvGvMRz3jKwTW
bLU364JDtu//O3yqE3OnvMk/aKZkQOjrf5F7ueY4ivSXFGZeP6PKqZXU32PaHrG0eP9OzSiIG8Gh
kvxXWyGiPL2/4OSdnlHMgd2sICY10ZlJdSBUA9rGxssnXYXcG6GsvVLbLf2tViIcN1Xggviukr1F
e6Su1IghbixWdQB+EN5iVfVhHEFZcO79Xn0X8R2ZB3GiCmyv6yrR9J+kh4B2U3UKbcbG8IMNMoFk
3Kc7U8sNwCqnuQ0XV0XnmbCWSvdbzxfikMf6b+hbOnv1Du5gel/ITNK05G6ihOqU50wRUWQscdIJ
jeIgUgtG7R2S/xNjo/GxuozCIyfStK+KHOQ/wL0UXiCCvpJQF6epHaJmOsT+agfe1ACxpajLAEfp
He1eV7rU7QRelqhLuIMGPrHaGRensZ6pY6aEJ9G/7H3cFEUcNPyQITf4PtuboVln7dH3uN4a1bxb
2M95KmWtKMeSS8/jHxTJmnLKLyV9KQM+D+hJX7Uu53UDvmua+aCh1xjTl4/tD//mcOiJr91g3et6
62mL6b4fcHHmcrSFVuJRZNIZ3oG8An3iVWT5GpExJtKiK6F7NRprWsJBSaf8EwFiMDBeGLvQjLyI
IlE+k75Iv0DsO4dlr+mcrfCLb/gOYSMK/1wgavRSHzNCZ9FgrpsaXNxMVmIyuD/sgl+5xhjb74nW
gHTgxNRp7C5EilarbalC2XwoDqreY/BoeM6x+aOW8wvFyGcMYImj06Km/WulJangwhJN6VwZeKZI
D4h4SdNvXnNcQHT4zD++umZhIORM4kXpkbLwp6+p/sY2hVsyxfUpZ/4cEqYhqG+jJwOthhwF8rzN
+Jb2iZHPc39lvU4ErhTK1K9MPbnmePnP5son4rS0R4z8IYjprotsyN5dkbV63Zh8CP9E5lozeDC4
1yOiQVzHJjUa32tjvnppRIOUhs+RDzZGmgH+4NpirkwJtkn2a62O+1klkZPiIS8blUQD7gws2uDc
Dju/M+vKtfMdWN8RQTTnUzlRitBOu4XBIJAxHsIarER+mUWx/yfxLokBN4UY9KOZs3AY2xMyocPI
sIZsRgR0f1CSdX+EWwaIz/4rZPmRnzjV0uBpjXUm/G1NojoG57hDsYQSQQeN3B8hlY9M/4+HPAN+
bxE8vhzNePB3KdX91aD3ZvJZorSbLhZyX2XFJk2HVDfedTJmbZpWZ/fMVBEwvQVPIn1SPqToxotk
rCE0giRLbv6papx0VFePAKsYQ/1rWCqlyi6qh2tOkjEVAO6FbdphivwUujgagWSMRtSdIdTYcTV9
Po1yOd6FYc/vq/5PPopOKGxU6KIimkIy/5CBdjSrPUzmcw7L+jCfpZ04FuLwavDeDX7CCPyokR+Q
zeyXqo5EXLBo20eXPiXacZZvpSk0isVaEhUIuqZ7NpRvnih88dP5CeYlgaLpB+YdlszgN4psq0UX
v4lx7pqciIQ7STWgOsYxGJSR4XXTpmsKg3nBTJYkEZGLIdWviuohTIKiBOKjEtwD/vYZV4rNvrYQ
Bnt4FFXkxvZyS2FE5qrtknOVrRbrnFi2lQODbx2i8riLAHmbagml3Eo8ShkeKdeKoErnPc14yCoh
iTPrtQpwaFf6vPVbiL+5JxITs6qdicCAqJz2VnctRumJlgYBK4OJsVafY7lopFYcboOvtZup7Ve0
CDc/Ht5uQ0Zbhc0gq0RI9wi4rl3SMPgYmuPsSfYZ03iyRrGj8yMdj7NylVUpALaRJaK7vTafpgMW
LQuY341dF8Qk23TkSwYTFjxV+JcSrnls0nXsOeNYWIJDDal6qakqiCK3Gz0C+OeW5b31cZtu2bQr
guzIznURGseEvM6M/eNzFcGasAJHIubWBCqhz/mkdjfR+mmcKVrYlbLuG2ok7DWz+8RiMXeEFO+c
UfYZS0/4eKKwln252jDVUVp0612eGIpQfYgPgFiL4Zx13AWGqoY4eJTcSHFx8neYAuDDVJI+KHxe
9kpeuvT6tWgCnDc3pibsrlkkkzfXqoGAAOqxwK6I1Kz83AndqMckrBhyUri8T3Af1aHylxUfoc8x
TERTMgCi/FU3+Njm/KOtdz5NqLCjk6w4QYMBJqjpthV2QOKgm8k4k15V6gAcelrrAaI2uYwla3ZF
I6yU7z0YtiB/dzeyVNm7jJLEJwvjYwetvu9rBPLlNmZpgLpeQY0YqG3P0ULD3puqRhoFFLw7g2FD
FNb8YRWvOQ/46K5aVIFh3x8464BriJLf6dP3fF/q75kS7XhtAlIq0CB09tpRVKcBScHLrAqKvGo3
J1nZcnyERMycMclxvsEb7oUMpZfTEYMj1IjsZoFkkKGS2tCMuxJv8QRYHOrtvO/+lpid7JBMkbjy
XSwc6Qvuq0l4xTv19WUb6ZFnaKKHaaQiknKc360i9hsSBIcFpxF+ylSJ2X515at6lj4iGiT2UL7F
O2wOMsSJIMA02HCFH43qD9vgBiBHjfcju8aXMT2rcMO5m9FK4a3ukwlT+Ez95f09voaHZvCacDF4
bQ0Wp77rAIhZDmKICLOP6kuNtLccpcuBpEArHNV/YG8j3F7u4oTLukxXBDlHkHLxl9QJISoXCo43
AZHdwpq3SZPgQ3LFznyPAluRjHf7nvK3nkC6N58vH+VNZCOX/jemXjgMsbmJ8gi3Tq/ec1Ib8ru4
DMKud15lN/7WZQozD6kKRd3rkpQqQL50MxhPVwJTorP7NKYNKp6MFrmCt9hurZRSdoVQalTsQmAW
Me3bche2hwK9Yp7DCGTTJXcCXqtlr3vcBb4PFSeX9OstivIL8C3cimSGg5U8Ws+f7PiglVjSn0he
k80rY4ZXJ/6JJOr8WmIS81qT4GitiSfVVPapEveLyj0sVdL+gr0V6/UZZwaOAkkqvqWgI2j9M+Sc
Tm4b96FDJ/3KTsO9rviYuPGdGkms+e+kVaRZjUps263R5plJFVYCsO32ahF7g+5so1mA5YIgDFEd
JyppHTPeOwOSekXlcdM9BGQVl7cCAoo6aDosP6K1SBk7loKSM3yvYJ4a7IVEJIi9VmhKI53UZJ48
fsUHeo3n9lwZs5Wsom8w0br//KYfDQ1T0RyhzlKrnxCoA589s81BD4zumxIapIx7ttAk4Sj7iYok
vS94VCdpEGaWrlUxiRuWapFWQ+1O7XJwzA5toeMzeOyhAJ5Uv71I0PXBkGUgZNxpChMbJp58Pxdv
GDCO1LMCXvGKjcRhuUIHg1KZRx3yl/wIFNTfiBme/bX4fSyA+FIQelaL2nLx3diYDfCkmEmTInkk
3Tt6uL27srHvFfvFIXp3Yr//WzPL1GVxtwqUVYiQSRR0FzQg5FxOBRQxHZ90KRQeGRKmAQTVcTeJ
qXJv3bmiPnw4nHxusa8qCCJOFwVgoXpO8uqWclQnNyfwbWLwkv8gq+a7Ppzwhk/Gb2+vmQy1g0rP
Ou6cU/+TfQ1tyzk9lihLK43hbeUor2bhegmuL5pGLlDElAwopx2VRanoSWUVtu4phamp+64OA9TG
uTz/eSV1rGQFtBvFLfMGxhrWO4zYgYnAgpfG1WphBETbXm8oitM7fvGuH8gLDKjmhDIT8wbMiJWw
GVXTDqqAYgMRdn08zlZIWmO0bKxJKkv4OwFjQTt/9vm8nLutR0iBlQeEDPSeDgPL8B2j/20U5sqE
+kCGPo8yqa/uITMEceAylIAvsUEZIETOycFSbKwl4VvVNqMJD1FDSd+29cPDiyxFUZXc/8MBBuaW
St14ANYpUPBenT4K27JRS+ockcekvjW34DYby2EnO0oC0Am5Iz9i+zSbAgXrz0Az4CpOfCuPc+1F
VEI+WBxusZQ/uv/iwekCgwcW2rUlIetsKHb8Cb01BnTyYjiUcR+7LSSW8og54eJqTtd3tk/bDFIz
qnFuuDt+PeZZ2QZv/b9vKDPqoS5vleR4QFVFagvLSjMTdWtbO2lrCTYGVQIGl8taYJWb3Vqpcb24
7r1rm+IkQoPPgt2cSgg59YdZu/NbN3vi6S6RtatJT9D47mDBCnb0ZwEZT+wU1a3RjyoiBD7yCbtW
IUeW30vpW7nXKlq1Y+LTlSREvERN43JhcASebromTCSQtiOfBALsYqfQpXArCIR0BLMo/ZS8UFP/
toJLTTNRHYEZWCZHemZyiCFz5J7FbPUq5YFJkpBB8ItAawNf4ZcZ2ZtW8mxVaQbSNDgzlvW7TVMd
wjxWrx6wRftJwtE3tfb6+uU+UZdY8Za3Gfy5cnbDG+JQOWq503XyIon85fueb6hQ+MucYFAR8rMH
gtc86llpIJpkt0XnAqSjq97gTraKEMjj6FPso4SqUt0+YUoiekjHLw6zZlZRnsJFo8uKx4BePB2O
x8PS+f6dbOhU3/fHTZBYn4Q3KozlyZSmv7xuwV0S/erN3ZLysO0PLoiWea8nscf2IITInjR0ko17
9qaQbaUMLSp/Kzs7NKIAHK+mZrMmg2gJl6/CG5+8hUKPBfvo1clYvBM8l3CZSA1b6F+xa/hiiHxb
q6RVvMIRDXSpNXrYB7pfkCwY8rCsoVX+B6iRghb6HS5AgZiwYxPq3qKF61teP1R2Cb65kT2YwrhM
+pSU0+xqHWAJ3tdnrz1KJMiJ5WonO4m5uwkTSonAsUdT10SQG7Fx8MNI/IOly+MD3ne7BapKteX2
NsHHex7KYkZ/C6k9vfjbfCmc0DkTmnkV8tkELBU5iXlphDQmbALJ4eXeI13wz9fk85WF4Er+XgMs
GObQkWIDpiCc+0HSgKDSATasZYMmTCLKrm2ANxprNW2cnDvNQ3VROfdK23FezqQG9BA13S0clOVh
x70s5DS3lXChcmS7ceUBk6JbcIPdo7hp4YrVw2sKM1hV8gQ+QJI7di5gvqrIW/2ES/5S0X6MyIZZ
XUeevGC2KMlJ6aV2ZW9/XE5BEl04A8hBPHvtbEkkL1D5bnd6qYkYZMn/zTSCD4QJEgAtSg7yjEHl
J2IVeO9b9dXW0BJ8QjWiKLVCXYcVT3VYPt3jJNFDYTrQAHZB9Jt+6coBOCfuSF310aojBM2bMAVP
WdxiV35IrxWvnDoUBD6tm/lYCKsC8XdvEYbXrP9IE+5399OYrFjRis9yDS6S8GS2fFjzaMcIGKQ6
/4TJKP0bq/QHQwE4spBbnYj9ae02sItp2g5vBQw1U57+VeYw8gvt2ANr3BG4vNGdB0uB39Dgs7cY
7IS8FqkGKM13xw51+fBM/LZtENqmfye6st5E4y0ZX7tG8qXXPhz2ZVGzlDdQInJYkzTyTKOMXe39
VTX7PFbjK4wr+C+egaVeUFm/sTgeHKSSi0vaDmexoBMMTFVhExsflNz+QEs4zscEYFaWVOW/r1NW
IOzTvXoqcL11rudwoy6HTNrhakD/PJDnba4bNl1lClJ9yxRBq8lxnHcg0FN4vMNXRVZVi04d6Xph
yjKXab70xeOn0Nzu32r76hcpDeT2njQKy1aLpRBW0hv+4urr4hcYLREO0fAAEzAgTlA53BH+bdUo
mzckAxlFKg1Y4A1UcWbCALYyehlX6CljIN7sTIRjUFhyosJRdqajw+8WJb6gWkGljzgwxrG8fn3q
LdKF5K5xjhQavpc3s50buDRo0Gg5YQmaJdPhrT6Vq4VuLgT2RVmDJecegs8zMiAAg0MCe1rqIAdW
wL3ZT4GPq/gT6XC9df1bXNmlyUAk+wXtLpF+5LckKJcTP1PhrnrCIPacN/6Exhaa/XNjp1Ud3glR
fPyToKA04A6PFETO4XyGH/FJbt63bq4vN737Etzxmp8do0ULPCqsaV49KBaT6JUKFG693qppcizx
H/zIipeNU8OUra8bl3ec0dY+a22OnsBKvKthcOEQcCszYKEnZvg/bXYPgUbhDwe8c6XvfkgOHijp
xDB/hhv3CeQEdNcZF1u/6oynvjMfVTAfsM0h0KIbBxDYOSrWOSSl7wasyrGggspQ4/Agdq6eKogl
OkHRfmSnPs+SnYm0rrLWDbNI3gkambJznVIQR61tRPypmg/kEX+diPOt9N1gEyNA3OdJEpYt/ffW
3UvlS8dlcdEQrO9M/fJB7WqN7RXENvzWpA+D3rf6YfVlBGIHpTq2PDKrwhfQ4SuL/MhMiSJf8QU8
yfTj303BbShUlQO3q7TjYE7ylA9IrJtJG9GU298WsT6n3yGbzpGimar/S6kitdloZECM2hxi7hqA
sT4zFnj2tK8E65qj6Q/HIm27IeG3GO/gg1Q6cLNW5Fb3liETFwNl50LML3i4FqRgfuaawlkO20tR
+qaQqOV1aFl9Eo5ZKuz9XmC+krs6CTqkrdAVZafem7qul8jx5rLbqmv/GVEsIyAtWbOiYJ13X/iM
gJitbKdu2aUfCguetHBbZtOiptZKNR2ZllasYMsR5qTK/79EUosChT93XyKRkU8WFn5NdH8XSMWR
fpud0sgFwaxGR42EqHzvlcwmpaqytoLaVttW4Sp68vjVhUfqEWRoP+ziKuxv/Em4pZABAyZzTFWg
3ne/ssJ/kst6bnkKNnchdohvtGe9nMyKz3nIUsgLsBRwtls9YTHADdGLRkazWTlWMQVE9QffzUXf
QdoFlRd5Z/hzsRRTl5xAyVdYj9RrZ4MKtqYmo1ntpH/33ahOWJow/P0agE0MVqn6VYViK8582ybt
eAPPI6c4oQXhUc9EoKdEcpz7CdaBFrJVu9kcxaM8VxhUMIqhZdyoLMJdgQdKBIWd0FXWzEx/HvfW
t9DnyJF9HFZJ/9vOOriWwQ4jw6wFyHPeqVA8SFYLhWgTqoTfW9WXvzJeOs+EGZrzbIbmNVVtkfQp
Z3xfnq7tbjaBzVmfn7PKkjI3C9Tv96LKgil8WXzJoEK2LfBHDnLFlj5eGf7Dw/UUzQ3MjLk3Ava7
3ciLR8iDzSP8HuUmYwsN1FkHs2iDALkiA49loOaC3kU85XnK8r0K0ui64V+X54E+ligWq/nyCk4+
W6IRhZ9c/I/oBSDeoNiPhY7RyL4WuIgcJQwvWifpSlJQl+iRxOu2a3hjbIXszpn8lfmoyLa0E/mP
z/BdKdsxAisIDWB3MuGBocEvWmNBkryylaP36TO9Ir6kzHuhnhk2MdGKEG7Ls7ARUT/P92cRQB3U
zOarKm0T8uF9zUR5usqRQwSssu5Lq9EGIM4W6RA9+hmR2Oshpi9r2/b9xQjJUlYR/GZU8V88n3Tx
pRpAdSgmW4HML3XpsqektbbVGse64rJ+RmyRXITXpDQVnE5Wumg03aguKeXdfTw3aYDJMJT4RVlb
+iPGNKPTBnexBXtXKaJaGkoBXYe99lgvikQT2KubjFn5GxeCwnjXbRVxlaZXBnHF9cC4KaTF8K1V
wdYm+FhRwb4k2dPcKa91AkGmwVORbRYp5zBkFcPClbM4xSe/lAmKql2yUkeQIoq1LvgSSvi6Hjtd
Sif8nZMGnK3GsHwVOVqHiFJMWgxP+Ii+nU+tuh1kqYckjOYuzU/YIWON9YUlGaxpm5qk7i581lJA
fItvuE47CjeaUsRpP5AQQ0R4C5rfxcRyJpbjPngo70yON45nuIH7oYsJkAt0H2hY/Gb3cR2skQqb
YuBfKBHYFLFBKyZ05z+9xuudZZOsRhqrJ5rhC1f8iNmAQrqXgOiACP8xuX4rSXBOHPE5iBSqlR9T
LyhaPKUaWtwqZ7TDGJqi1QFz0UQ//nVuJ9PqZ55DaY4HWbVN7FC5dm33ascl8Qd4U6oOWDSoEand
lLApUPcyd/eAowklFqhpl/oR1j3cy9ZwuzzgAHwpy0mv0C7eY9Qzr3/53ROkY4nie0R6c+2qx5+b
W/upIgfTx/40HgBR/vedPBwsYWH7+Z7q8W+ofjfJmCNxN0KbAGYVpxb/J6u+SoLKu5dzF3jKDo9J
WC2SweKxe6JAL+ILZEsPWznuHlPDq5tf5w6e3qcnMO5qspUJluqM8kGJloQPkkGSMUO50pAZ3FzX
hBu4dND0r3iL0JlXzm9++1c+9et3kYJv8XC8/ruZj9YNAYZHHUy3dpQ3KBQvRbOVsdi3zYK8FZQe
D5eka6nPFJAfLfEW86rU1l5VB+TK4XKY+n6xy+mlI24nYbgWMgc5c26de/lbkne/kqYfnuEjtjAO
k2EtcNxV6MSPW/0X5jL4UELFxyK3AR4Z9h5/X2yb61yZPLHPlTj6bUZAlidcizFPTyn2CHwvxOGN
0HBtZdkbsILDnGtocMYJHDje5rXKUeJ3GlIDuWeH2spx0e4rgCtGUfPQXSggcGnmQEE2NMxEsZVu
02102ErB7vzm7WrKk5Z2VnLFg2bYDu/QKnyYR4c0kCa908GCpG5cN/gmndL3SIXVHJvl4OGvNCxq
MldkKqhjLyJoE08G3Rn7jbqwZiUMtLdvs8v3hmMQoqwBh4dhnNevGgrU6zm84DQ9Ie8N55iWIZCW
vWrID+SN/rxMcMVKHHIXUCm3avb3IMx8K6kK9b7Do++k0ED7jFJ8pPfD9OWB0a5Jwc8ZXixIBUp1
SShl8w1lts8WuGUDPxuCMkoNZpXS0rjhRiFrH4hlaqnv2SV8a5HmEHtC/Hxn+hzaFLpGIgOrIsIU
wiKQA9UA0WMvNHb7BOSYO041sH8Ag0t0FUzJ1+tdCNyYJtuzcxY0BoRd85jxxi6/sKQHuXJIUVi4
6DS85ofULM+HRZSLdVFP1nmsghusZMOmqKWcA3J+on+0bv3T2nJM+rOk5qpTzSOCfwaYEDkhSTv5
pmIeYIKZgOFiO0c7sfZ2J5ykPG33TIrjmM09o4/3tsmUOmwn2x6Z5WiodGWDO9LA28ejjP2lWJ2e
4WnGEUlTcxfNrLtdy+48jvPfo7vWlcY0CcMCDRnKI5XhlNBfAgsNZSVw8nla+pN8hzY26Gqtwlpn
f+Gm9xlcvyrZ+JWWvMddpKVPbu65MCA7FldvCRzks0aQWtw8xilG0QxHPzlm/ks/lN4YJjQ1vwHH
6iNb2Fr0LZ6THy+t4uX2CofW39UgP0y2q5TB1trgXslLtJvRyGdhk9rlLcC7PR0qJPBn8RsScUki
A6TCDJJdY4Ksd5g+7knLbCztKLeEWJ2TU05yNVicifWQTIYErwpnbgj+eaYt53Ok6nG0Lxvb4ls9
/ccwBnFk5iBLYyNoSBOOUixJfs2i1U9/7sCSOwtoJupnPXwujMxQUKGI4HTxHOoC6roNb85IuRRk
pNRaWjCGn+9eq6GvB085pWlV6xqRZfT0E3BjYIuXmjSPgeiDNxW8q3PXHSLxypFI4aZDLgCU5AiI
mtF7NxxfLL0mCs3PsEBL2bhbNEo0Mzf5FVizocMv8S5K0gal+5b+WNWAmnYY+VeATPLr7yKmjVf1
0ETprdBR2/Id6RobiDNGk+JvgcoXie6GxxdJpWrJcomaDLqadGTHp/tt/E0fMJqUDYXCTgYS94bS
9Bp3nB8J9pKfIvcOCLc6YnrdJT5c9JOnwlF505/XSQVuasPcyAb8LfnoVm/3ieD93BbFo76B6T8I
4Id0HYiw1993llqdp/9be3fXh7mAUJu6TUjE4mQQwfpvQn520hiS0HntgEIWYekaKsbdLxnFa8IK
Lxkf3KS3dR4/TjHyADTPivtrDzn/iQo+lOIfwsasBKNW+S9AtxYJoKXTTDj/PEX5GFTec1IQlaDG
S5+//FOzifIn7ah3VvbeyrGp7B68chRyroua26HsgForwwSdTN6Avv0ai9B7tIhi9v6l4DIf1HV4
Fj7TzINvmbHltBkhhNLBoyyT232eSUu8iOgwgIeN8lNvaRpUdeD+D4hsagGUh8TMfeKswTC/8LmF
rt0sFpcK1ajdF8p3vukb29PQqSozOP7qupF/D/kBiJuJ4VJBhC8NguyEwvdOm5F74sgYzJ7eDf6A
1wSY4jVbTB6IjzfbthYZWN0Lu7tRx9iNMfeLx0x7AbYkJIBQI0uuFyv6ib7sc8mbm6WUlbQylMvO
XLhk+4pYsn+nrT5xgwNuyxtanzQg89hGh1Lv8sLndSJ1xA4xOfTCViWsFgYbOGZNfgnoz/kuH4Wc
tVgIyMc9M1pBj3g4X/CdBajuWPMzu9KVKtZe4GnMbahXILoIIOnaFUxMYaPBy+SvlKfNyTnGLjLD
+M5vaZZQi5bIuPsPsHpcirzZRTL1qqvhAQpFtBHDuu7sRrpDzjLNi0gMaJCS636h9TvA7gZlFHFB
i59KajqKkdK31MP/h34oNZ1lbpBcEANKOdkcPDWkdujaWbFIA8rVe9qf5uS2WoAspxpyCnyGA8Ct
63EwPZBi87Ngko1ElR2dQUHVuLHHpnGr66bRAZ3CxvSqEY5oXB1j5z4b+swQ037XXUs++JGDExiE
/N/OQPjqlj6R1eHns3l3dnQHbOcEEft39kRXcWxQaSsRkBN7zB3kIt+4irHwijr5JKFJGMTn5nvH
gFMbq0Xy1SR3aSNUWF/7OQmvu7ojvMMsEwSFg2mkwS4uD2WbTl34ucbm3cgSd9g1WIlbCKCpiIbc
JC1gwuG81poFMxGkRvbkBrtiE221/XFhERpdS8nKFndoXSKVHr9mbmLyxsgCsGv5biqfl73ThJU6
+Ih4Brv6BGjUzuqexnX4/L71pbn3zOWkoidCDt058nsUmqSDXUTxiXU9fqe84LukSZgBXvmg23vH
LCfzQ4fSFFLugLgyWROuemX1rOWhyrBnnn7ZAQZXvvy1JGnj9ZVTWlTE4yyrXdWWQPxeiGyRt8BJ
AB+j2Ff9BzzwyTjDTuSpaQ9dzekmWhr9x3CJtdv4Nu0+BLEOkcRWgBQKI4Tdp1klbi3iMbTf2QsJ
tgW5uMjAR2Ag3h2XmjJPM4/3il4uhC0XAVqLlP56Ou8ZJHVcUKAa1+rReJwSd8zLNbQfN+byqjgo
TCaMNN5bxfJoxJGCoPaNa21P4VszrSPN86r/a2fSzSLrAb3uQshtphCBZVYp3fHRboNcKq0ph6VO
cuW3KPDj2sU4bniMwsa18+f4hbjPoevJj8IcZsK8Pk062M1mW8Sxx97yGHQ3LvFg6/wlX+6GYfLH
Gu6kTpf3xVbSrqxxPu+GBsRMXx7Cut/s+1CFADeMtwhit/fIQ9cDeBd2adCxGJKXbqQu+IJWVCL8
eAmyI+hwVe7rYvBkLhOEWtvtcPfpY8yHoNiMMYWeOlXTdpzBPCsXSrCn3wEn4QxGuIIAVJdO/jrc
4w4ASV10PbK+aQtchRsBSOpPgNvsYB0TkCAS1jP2Ynrq5jBa/zJvRxVbmtE1Um1OsJOI4KTw4Jdg
6SOdfUXdKHwUHOGY8Y1qJAy3P1TuDsk+jSQLoR98uzC+Ul3AcEzSDQbOfwgrxQMSjtVpvKrC0rSB
4alEFGY4emn+JhEZQL4i08nBEFjmbH0Gur6Phw5WXl4YRN0+6kwiQzx9H43mbLI5CeML1BHxe2fv
2+TE06j9gimeJIJfJxlOhc3ytMtHwhCcSQVsKugHShC96IMasB/38vBUGsAt1Ykjdh0XZztqJ1X4
i4OsUh8QCnWTEtlNh43Ltd8w3rEE+LXfC1nStXH4WAsNBd5Yh0AkFnBbLsdXd+sPfTrh98jCxv0K
s/0K2gCS+ZRC+kHu8lE1eOYh/56Dnk2Do5/ZmE9ZuZZDeilZFj5kOzkabtkqDJ5RWVVf+HXyT73Q
66JP2unWTRL4WstIFd6S2qe+A7fgDVJrZoEhit6wID9jh+rcIWAOPnMzLQAoQ1adszBGnDFRbLj5
ZxN8mlgNAKeYvorTHhU88qyv6KTnBs0tWnJb9bd3gAohzk3cWutO4iqfI73Qh0vMHS7gApqxeh8U
aIAOH+e5t7118BSIqRHCvZCRgmHF36eEx3EyKw2FUj3FpCpxyuWY5iMMBpacQHNY92kZcTA5kehI
Mzf8wAv0IagnBtay5JYsccZyECZ4cEPVruElkBFyFCXda9a9hgHm3WyQtbGmjhFIDvOFCvq9PL/a
cDKbtnXLueR0lucKEnYTFEWDwdWozOl4UakzqXQHNLJYIHL0KDiCEvKZf2C5xyekStUOT7ZqwT7W
uJapPHyfDBwg5UCBrENKq/bubx9yKMvNcfJK9KpzGn6VF3B8bim9j6wpultpybi45Kj9jGGp4O63
eGElap40Y964rcjkMkJ0NYeadNXY2cq5aZKQxHrYBd7G2Ljlg1p2BaxXVxXLKYqYEbCWIZq0YZYT
864wWcV1X/vaOJu9VfwhWcWu2gaJu+ynbVUhLFWb1uf1saf7gefH0rbkSCPvSjmFPr+6a9H9WBEJ
6egj0JDwkIict1yDEOWQ+X4P1zxui92uK/pT2vfgLPwA26gs7GxUCLlzAU6jm96gvxfHze4PxLBl
W/LScUr75bjtNIMOA+0XViqhf0t0qE3/v3dqUjHQqi+Bb36HGxjwVwJqNT56uMM10yIGVvh7acon
DScFosgQDcxCYoE8W4/DVYLoO4WLKgEszQ9f7SsEHWuzR6a9dJT2+o98mcOnGOu6Quwx5uDbDvbo
CCWPK6fQCAYN8ihfDCJX6/x56VOxlNLtiE4bqNLGhjgLjeii0NLVmqBthOxyyo/yZMh+AJPTskd/
FQjL52RsqtcJyX65p7dCJ5SsPAFRErV2yybF6dMvreUee4IyO/tJ2cMGI0KbyCvyXY7CROwsWlzL
fPRifti45gu/iisTrNwweh2mqi7WXdRazI4zDFqA0zsS9AkrCTZKWlqrQITa1ZDc32JlKpir2R7O
FfdIpnh7FNp8FQo3cRXcG30VWVBG+OdxTej2bkMyPSWq31q+LqdoZCKz9OTpnpkQT97p8V9z+Hs2
5rnD7AI5Y8uoF07ViDxJFgMcCD0h3ZLv0NxU4ARTIiVweDEbG0yv3AgDpt0MZ5eWnMLrl9D0rwkk
Yj8R45SRee1R80eMXMrPa/OiQX4b8z6nGpqbQJfWjHxAOylY9n4+cCOLMcrBm30UkMmK4SWU+5d4
QhN0fx/jt8IyTGBXVnHF5VZ3ouamInLJN0zRf0Ju1TIR0Y//zHXzY+mDEyQWOAllSbWxtpRHId4N
Q1J7bNBlvgoCBJ1MPML95FXVsb2drcOEXHU4RSA7zqBlPpgOcXd6jcF/U7COIru6la3h7O5h8zdl
CHJ/8Gjx4fCoVOZcDB6dFN+l+vHv8yACTIKwsQ91TYSGVbM1DYznnVwhDDjU/qJCheHgZjbW2KRH
9Mlsz8ua51zlZn/if9ROSI8Wz3TnOPPxo4Ql2hPQjXpHPHsSrJQWRmwVC9XTF6rRTocRefLAgtXs
juvxNmjEru0ZqOjSIzLwRHkORpjUsl9RfJ9MRpw2PdUlrXyGa1fjjDaOSzwG3wnVP+1jnFo+XGoB
vWA93xv7+0o5yCme7aRhZMHrFWrd7N1Pmuw36OVyF7VGF4hx5yC8SZuK3xTxfM+DW80+vhyiY4uQ
v+FlLmRBvmTn01ADhoQGgAOhyUziJnP6zQe2GL1ubhS4gGpDJeDfHW6r00XTkkXNCnqOc7zJYMZq
bGPEDFU2Kik0rkF3zEC+N2jJ33MzmwtVGfBH6O3r1mV6sj77kV8QHbYw9Nk8qUwf34nBQSIp56Tf
2h4k8PuyfbrAY9zwA/CGLVwj6u4LU7No9GLDwNLwx4fF6xzd62xEsYO2kLJV+3HvImtn7rG+49Wm
c/vFOMwRz23NJ+dffRRfKZZlOmnYtL4Cgonk54/cUGvwd/fDGFvVFJJC+pxeH1UeK8SuarxFCl6e
tLRfVxa+vdIPql5T5OYtBJM1N90pfEbeoEFdkp+h0Wf69lA8BEF2FC7MukfNpeH3EoX4d6A/jOtK
ttLLt4oIwIekM0R6b0c5RD76g5XA5vYGxUSzaz6NzTfOlk6sCKZtaTaygdFk985KrSn2l2+LBYnT
Fx6BJsvf2GLF/0dSJXSVx+YzGZLCG/9nMsN/0kOKCQP+UjdcvuXFj/bxaa3b6g9h4JkyRr3nFet+
n65uhLrbnJr+k2wC8t2V/nUp+9j1c2d7LS2V0jxX4MsGuYiil7cCyaAguay8HVINpMRB+74Rrvku
cnhgLycBHmKr5rLO51EkIMryAVzOeZLXpgSEZ1nwMablu8CRsDRBhwuKxj249vLvWCkWtLo+IdXq
oWVIksLH6p5fvMLQF1MMnh7sqBoC6b2MdRoIFJGBgDau6InPNpHYsPvD0KzTXzr+bFYtF9SwaXKk
ycOGxfS5gSEjtVvx0Ww5dzqTBqe+Zml/tsOA7hKHGP7HiTJfbkD/AdT7teQlKopAsqopDA0N5cZL
eLXoBfy5qwFYM+fesPdITl2mOAZXbbGUKCRcsluQran81lnKacw++PeYQXnPFDj2yPjfTOXBxQt7
XlLCZ6QwN0RQ2YtAOhV/URDsZ6dQd1mbm3KtwJiOqn+k03hG/HlIypjFCvUCEFnqnOlCmlW9axcu
yUhz+J6HNCWVa4esI6AYqYBnRTq1ic+5Vbf70fr99J41Pj9AbLcaCC0yFZKOXS0f/kPrkMG5PUeY
ZiGIEKEF7MV7RKZYWhGSvW0s67Ur4E5tMjHcLiG8ZvUl1JSqNaFUVU8LaBTgDWbDXguf24SDzKYC
xkplib0l3mDkeGaccFGwRLLMChRCOjs9sXbeZ93MOMzAjbhtfrj0fReMOXAej8WcxzmldyhgBLaJ
ZzlWhA72zlHKAfTYr1FUku7cCOwtPO1gDkze9IDQITtCwOd2lf5/ZG0RI7QsnkqG4FTGenE2q3if
kHr5tHgO616Oqa+WIgb/MwBOAy6550HBZz1L4LWv22qd2Uz0A1kv29Dkx4wjN9AaNsSRhidkuGqh
abNhm268Fol4HGTIl0ZawA8+4XAls+wW+uKTCaGgm7iKav0JOFAEcCWRRhWqMUeaRiodI4PUM2uT
NfR7CmWhFrMsS2Tjerqw/n5F/EwwPjX0r7YBJFISxTebY7959V2TvjoMrqqRsdefi5j02o+nMH4f
yUQQTykbBZ/mdLmNdWW+nAjOrxgHOVVi5tR5SQ8bIn4t6vIkS2swsVkXdOMgDhouVxOemY9CwRkx
oCyxJBvg1CufoEbsIDQYg5AUTxKwh2wAcYFjUi1NI7aCg3arZiwf0RNlvugH9rhOOfEUFT2mRqQW
BWtRF+ZioUluyvfhFNkIW5mRLPmC8FOh9+lOyuzNGVnrU/j2tXepWQA4u1fpubxKhuYaMrP40dOw
MKdqr9pfUBivYjRllg1GCkddAZYmz77wUQ9seDnX1jsh9YXVYC9iWFnIKke6EgEnRptHjvueg0IB
bB7nftg8UFTntU/qGtn3br6f27u5nWbT4yW35VVbp4y17KP0S7UIqjyg6/SS3S2uh+Az0+puUsTe
zyNEZYEEKVhPsO8yjEJBqfEWeZ0vFDHcK3+oMEATZkh18qlWYuqw3LpmyMxV5CM32xThw0teRuP5
w0nDEQR8CRQzEOjeqdjGkcWhxJzxweo1wA4KGEJ3EC8h5uzbMayYg+sG5aKin0e6hEQKpo20fLNb
17hB2niM7K6N0PPa0cdv2hZSm+bgqrHLbjktcu40riY9icJlKG8DGhm0PxNB2bVbZ/Wjmo5wB5T/
4orR1mN9NeSs5wtr9OOeiwjEXJyeXpJfYOrT73FgIaj4fFdYTCO7Ac6pkoqU/Z6R6dc4TRzXjouh
fFSwHlvidkJhIjRhxJcVN8UsTDhfOA1XqzXFyXAfrJVjjkhyoXm9Ioy4lAFXGXzvLy1VbaXnoFqX
Vsk5G+fNRiosS9EZwsj1FEJyRoKDvUpNxaICMzzMTZREDWgEnJjoFT5gQBkYtNxGVvMc63nCmRqJ
VpuJuHM5zHQTAT9HbrW1qgwoE8PPCe+CremD3XBvndFAhkh2Ex2m7HIzEn8PN+rwlP9rObf+lg+v
+U5ArsF9S7mqNck6l6W5WJUnlIqqXJtCO4VBDpk2yCaXuxDVcoxGzsPzFZNJzNUykNnwEXoR+NtM
j8XzYe+FupoV7DjkHUO9I45tN9GIMwn2EY4lvKnWx5ZZcPOFiLsKZI0kX1nbxJ7HZkNg1jYc/Cus
CSNSyA8UyofZ9k8P9+mrAT6DRZWQBIbiaM4PP7OcpQ6u8D7LHfaVMWnfQ/rpQsY5gxXPRetEUSBq
0FaxzqkrCFExWb2gDTOaOQxSHH/gCqJAqTZU8yv24Mml5O1FAJdno5dQo4u45NsdJr/hXxFae/4/
XiEUelML7H+8TUeSPc2QVakLH0/FFDa1veUYZxwgtic0rYIaY60ucO6LVEBK9Oo+BJILGS3a1jNe
N3bUNKyTC9Jvnwnt0vc4jtd7lmew985AMxlexzaE9/DGA8Sx5dvRt00d9h70JrtOQU0ij+3h0WH8
nRiXiz1jZyQjh11KdF8VGmNcq5c53eKZCBEEauMXC7sHX6FXWDazNfHiG/+faYnp319czZAHPm4z
oQ1aSx1fglistEC7Ai1ctU4PqDM1q9QeJk34PSF5YOEISjys0B4ljglXJDsDDiQCwkzB1eL93ky8
dVBrOqQ3sGjs3VDod1Ss0LadJfid09B8lZKgdCrGx+3cZ5ko8HLKMjWk6FT+qgWB30Kch3g0vlgA
G2RmfzZ5aTdFyh4k+ZYI1ELcRN2txVO5ck6CX84pK8mZVH6WQMFFeKIbaFIU2opemMfIFuXbji/H
sNigaH7UN4EKjW73Bn58rS2Zpnll07UsiWjCOKp38fgsPJPzHo8a6qin41RetU3wBrJsHcIMWbAS
JBIF7Snan48GlKTfu4QIIa7yVLJJ2WypzCwowB66GOt59AaQvHFM0e+ZJwgCBSG2aIoTqLGVH8P0
cR6chaIIQ0XU1RCwDWIOKU6h3esmDHcCNaF788aCsi+yz+LRGRLHdjxzL//WEv1a++gt1mtVYbXh
DB+kuCv2SuxqoSkD+rdUur7FJRb08IJ4xK2F0o2GdMCHlKKg7vMCWm7R5auq9LENhBlKv4Gact1g
KKho1ji+Or1h2zSdznmEVRO3wu1tFL/9h65hKUGWni2u6PAw/lix0aMcaHEgsvXIkzINRdTnts4j
TL+jmtbhDG8WTYVJBriHkMiZUmeNTJbvr2oGuZBrO7a8A6lI3NCUiSITId5osVUy+vuTvYSzIrXX
RRgQLUihJsnu1KH31pbO+oS+cjzInbM3/csozrmyWquj2Wa7tK04Gspp45dyBcn5kL6mt9C/2MKU
5iBCd99KzIawdfHFnjGPxOh2ZpsvR4u4oajqB0Xf9M55CcxCh5FBpAiFFl+Cmjvl5iRHcNSMuiwM
WAFSgL1pQqp4Y7GYSF9/6BEGQ6orpZBEeP8tmSNFuaJ7D7rrsyTPEFxBu7LCfPYDCa9YsZFh/B5v
8NTsek3aYJWW7P90FzwdWQBBqWa4cImrdgWAmhB+ZyAgr0dbByK/aFde5WNBPpuKHiXQToBhR4ki
EMPt54pb0W+GxJWRtRg6J08mGKmsql3gn9arqVgR10TVl2WB/j9qktrYV1DL47FnHgumTjKGvIKE
b75e28Bi2mohGbo5pL1a8GEXsjOjjnvNLrxU1NijhAT9Xxb74goVpbqjWW53HJYIrZos9TKXSJXz
3e6H0lwTtpHqcrZMedZ9kTdve62Usbq6iSfTT1cVX652QdnExUJGTPeLlzUytCe5RvGnrWdq0tCS
81ugKLF8zyEk9KFpA82B5TrNMmgBx3zVKhdsNPcuycowMvM1cerd2vmUaz+L6Jzd1lsJ+hijrLBX
M5D3PTTfn1rEqfmadEW3Nkljn2YhzsNEhlMHofebIhdvzRUEGGmFZxmvC4Qzjv9ivzCbmX+vMLgr
ODRsjDDucpXNCd8FONh2KNdZtXI8cotx/hTn3O2MVWoCVNnRlNKAbUWchlf+tKj1ljcuoOEVdUZo
byfrq5uJv4OaxJi+wPS8t59i9S8zdw+2Qx4gdPfRCe+ofNtfDMiiy8qbtAXTwHvj/Z/LPxwm9Xeb
J/EVuXs6kofn4Z/kdrXNQoLDTHD7oKm7y8atKv+MHhaowgmNecpKw0DBFXCN7eIe0apb2I0EJKS0
h2hXpgriEGVrYquzDSn5CGqDal27Xx1XQ28lmZMFyPPEVNG9BWR0D0sFTaV+RUi7KcfLGL64Pif0
i5bkBgf9qvF+BVRtZUxxeFG22+4AeNrLCnG+G+WULoKfyeYWnvqZrVAqOSnjcZvrErbsDt30TYgy
RL/KARkGhJrYDfHGxXUP4dqnfr2VmJdbmUpVp7lFGcvLr1scRzJnJR2ce8OO9pv3Avk1JdshDtBb
uWbs8tNCpwwUbQ1dm/zmkY3h0gm2Z5NB3wqutInyrGneqGkvWZ7GF7bAd2VQVF8Y1lAvqyubjj4a
SV8vhbSUQTpS/3Og4iQnRcNah3LA2HkVdOMel1RzRJ+P4aGUGeYaOLsvz1bcWpL2Z9y9I+3LaVYx
Ozh2fjAds9+oyUSfaI5qm6LkgKqW/P4sgyL/bso3DRC6Nhcb8EPAov7xZGZeOY7PjM2dY9QB3tGL
xmnp5pLdrSDjn1+t1mJr08xtP9zUJRDOJYAqcYo7VNbayObVx+YtU4D4CmA5E85dEmAKN8i+gdMy
4NTinOx1KbFTfaHvudiU98FcizFF9lzlJSlp0gRgOxJl/6exgXoY/BgrJa4Xx+0NORWu0Pdc+Sw8
jUsfg97aAIyjHBvarVnJZLJMYEcAojZ/fa4Fnw1dBNuEynmFeqvJK43V9D3HsBVri5vxyqpiREQQ
RK641tyLsZp9qT56JWARbZtbQxx1wl0rvZnlDBBqGpdCJ9cT5gTd0OxEsP9+wkrEclDaR3VNsyTK
m6JSa7WknpPrtbXqbFx18ys2G3nlK7Aj/3Kdeu4GpbVHz6P//2f9pny3RQAeGcwXHe48akP2+PFl
zKw1beXoGSA+ehTG5ejk+s4u0+wCsqY936DHZbeQeR3gS9UCNX/v3lMr/wDvKgL0TuSHHwipv4L8
8JYIzbTrRpu0Mqx7bEPuA6C7TdKHVHvkbXecs4/TxIlNy/cZSKXcviTXtBZJzrNQNgMle1mmG7nH
h4UL5nXOgby+6EdRzx1qnCOTa0xsTvhd/t62M3ofTOQGtGnFJ9LL5iJvmVY6QWBySn2CunMyFOGt
1jZBptiAgHPvFIiopYPni6Ike6pYblIhdjOKVn81rDQBG8LkDG2EKphKrG/uZ4LdIn4lO6JDNSx+
qA3yFCysrphv98CtLJ1qNjZNDmvn6UTBtc+QgdMXEsebsZ27TSkTZ5jbJPwz9GU5cMzJlZoHXwLJ
wTWX32am54f09M8gWyc4GPeYp69mB9arcLtUQdHmGWEnDF3UaJjdlYzxZ/57Qh39q7RDDDZJtga3
I4T0+/jKYHYi2AQshBNZfsFzFyUQ3rSB0tu35N5NUFFHjqS+iyQ9rLLF6D58X34NjUfEuiBHTds4
ryJvwwZr8EDirEXQgzX7KFnGO6bmu9i8go2uUeRnq3XqG9TAe+o77HxscWgiEkOH3XOXuFJUQoe/
QclirUkc3vBIMGu49uvNZLx2e1CFXNVoAtDV75iAdKoaqPGpus44R1zgTgFVFZjIoNIMmjAKpbtQ
oJ+AuYWxpLa8iL8bFXa0dSyQpszt9rNBYT834G/DW2nbAlzivu6bE7ul/+H349R3/0ro+RGxIXE9
mPRulVk92uD5F/PPxHXOQEhAx4suL8R5k2pYRVO6raf/g5qy22l1L6lpZGrw0G7GCNl2WWEEdrWS
sY9kI+p6C2Bfe7QspZmAPCehOUqaJ33G7ldC3E4tCKhD5lmz+51ttpRMVkB154UQ2ZbVuyWdIiOA
a14/lETFyGxPwe8tkmSTOBm3OHSNHS6dAD8X5b15gknlgNYWv44xc+nrumDEzBq652JAhzxJA5Il
msH4kBdO2Gv1prowUg0V22wFOypkZKGf2IXJNKd1fKm1VlcdoYq87L0Lb4PjlK8VUXM7OakH+nxg
CqyTzcUEZyGRamtR4xdhsPcnoOlL/07uuJvQS62SnTbSEsOINrVEqJwbHCB3v0QJ1FtygYDjc9do
3Vh7usG7gtqg4ECJo5kVyu4NccgXDMlmv/hrO27d5zF8023Yvab10s1D3EBt+7SIPOZ3H7mMEhTj
LOOtWjcGbOqzbJXyre5MBzYELsl4DG6BThjgL0lm6ivawnaOVgt9SxxdiYXHhWhRIoV3G00yzgDx
OxkybeaXOKvh3/EnTYU4LGxS45TulHxR315WzwzvtEK0vPxs/pUJE0+koSXBIy/Dg3GMbj8pBekQ
HYLWWX+hUQMp6lbRf88ORaEH4J3qQ5Co5zl2SBNUHtnXXpdsPRh6mlwCEc9g9BGMrkVrRHhi6oPM
KxgNAumWsDB8KdmI45bZBmyHpw7pXOVaAORo8mZ7yg4jTl0NN257oWH+TQrMiMlj1E1pbPHlaBy4
eUJIbX1sT2JtvOqAwvJ11BnDlT56bggWWmZH+db2HfNyL3yQ4wGRGLo04n6JiimPrjXZtwSodq1n
0Ry4nGySOCt+LoeFRnUIynwBO3q3nnasLHKq99SIB+ctYbXHO1tbPtQay4+K02LWKhgFHQgbDIxP
NqSdIfMjkWDJNqd1QDFBw+hOVMuc7bicrtTfFEBMtvcBJ4+V/060x2XmmIX2Ed9gZoEwyJ8MWkTK
HQvoOs2HasXrkQJFx1g8K7HyZef8Svxwk6mbso9vJw727FbLNnDd3u1zB1eXu06FPxiD1NDTFmQ8
L4TUi0B8YiWQmPjiNwrlsK11ytPa1FkMR16ngR6/J4rHswNVS3Nm78adYwq8ocrWn3BZ+0JJXqLS
tYtEIu0FmgotjmFYBEnEtr+laOrNzpwm8CNGErLWVaxxok2HM0NTtW4gsYfrT9rNG9rBJbvw60r0
cvw5RBdD7KiS/7oooPHwHdZmlonWhIr41BRjXJRCp8wHlR7cy9dkymAo7/enWc+k+KbqA5qVeZgS
ptG4/EbVc+xCOIFHPygM/v8eYf1f84vvUlNizlViAuYoWXpeqAkuOOiRo/Tes3UYRDatowhfBgqY
aKMUGzqf90z0uz66z8zQQl+hWez34iEWPzEAhTpNjMhvAxH8YWnJ2OGowd+YW7uZQiyiSPQJgPpo
B/v2EXYOocuyZ8vCWAyR2/JLIMY3SqmIVLe6TOPPuV9oBSLTj6PAJEhA4HIKnM7f1LYPPueJiLAF
Qu8w9tHXDhRBv5GE4BcZDU7/0r/MA6ox0HEePHyYvcXSXOlUic+UPQ5iflcnmobbRa8L4adz0/XC
RpF6CtGv6Rbs4/TGjUufmjVRDcKiYXP2FjYkH+xV+2lTSHIGPQIGmyTmDuiE0w5/TSnCpC+sNH5/
uy4Q3WJjnExzHWgfKTYKkkYaVHRgyfYDeFlbnQ5IyyFrjZl3IIAKeR4aC7rXc2gwth36Qae7zV1v
jazaB4U0NKA4Kbb16E9DPMcfBqFTwu+KPWgW5Ez2wHZFEzR6nwn1raCtRE+OIDLOaMQoaZ80cBIL
NyxDcimMW+ItoAG31nDhDJo3f2iU2X2JB8JbgTiBrhxjQtxvxQV6JZ1gngvTc7apax2LZnE7W/Io
olFsu64onIkwAMe/IRAuT8RUs2FcZKlIlYAvO/rqlckUNiozu5QiyVjFyRDKpM0Y6Ah0uCUVXbVN
6qqOWH6n0CczuC0lCIzpb7e4n6+9RFWchAcJLIdnM8ec4Vw25Klx1rtvZqPu2vHnj0rERXEht1Jd
ZQU1A5fmZPweD16vLz2M3sAFWA7sz3qTNmdqJDhvrEBjtwBUTuAHS/GA0vMmHAkHDctOZ06Mcc+Q
n7VRVtgTwgqXiMrWrUCfuoft4K62ZNqd5LHPdBhyWQm1IX+xaYTpnyRLeklVk1IRexvvsKcCrrL/
ddhQaLmAFKAoLy21QPqa+coDiPchPPQR4G+ZUYN9iTQDlAu4b8DCF9NQGh/vbP3cTCeDrqa+qlAL
f9VZo+saHAmQYNexyw/UNdFuLwZMPEfv+NVr7g5O1OQdiFYt8ppifRAb5oxHQG10Fq8q1v53YAJn
tNLtAWfekoOdoKZMinDv4goekTAYejVcg+KYW5rw0IgCu0rGUMHv0s5sYM4v5Ygq3/5TlTOXZ9Yz
eq+B7y0LoVEVSCPkgvhDqCp7ZSMxmc+3guqa5ZukF788mNFy9Fcbc/dTlXcZRps4RSW56Cw5amdh
P0Ki2KZ+T4HOx6OUPeNiG2R6kktQKfyCmfWq6UduP1E/HqqaUh7tWhjKln5P4EvcHKz4gPb2wDWS
oXLAP3RvOVX1gfgReGfqIjsKWm1r0+qEFtRu25QL5vK10wXbmrpOOf8LZVn7RcXuODgohG2TrJ1n
LSds7VfUEd2620GPTF7SMiPybFtM5VlVFALv32PS6Xrhl2/C1WdJuRv0J/Hi6ZZuHXohm7KhziNz
lM9X7hLgTFNmBLsphW3N4l0geLrMRNxKe1+BLqrGKdtDXV2MXOZnGqPKDqD5UYan0V56ansOtPcU
EPoqu9usDS1iDER2DiWOvQ+s1+OEvfiO7WVwYzcg9sE2Og7KMQ6OzGp2fGgbJtuBZeKKtyNXjVOB
e+XnzdTljmbuF92qKkjZFq0dwW4rTi45oyJs89LdE3zHuruxK7KOGhs0gWWcafq1fhvHYF0+NRnt
Qsq5wyFw5pBUjEIA0XX+1gb4QVYNBZRS6lJjyrVdheUo3oZR6hJpyK3kyyZ3mltqrXEJjygJ+KrT
1d+OtYtFt7pYUeOTWwTg0DF/YO/mLFK/qcArs0ZdAKIJ32erhsL5oODjt9l+JDztf7qM6/8BMr4U
vtWRkMfqM1Tfqs49IGN7H+GaI/rnPQTY/PBVEZJoGyOg4eAZwEXRRxflwJEvEe4rfaZEM9o8KNdK
apmKTrSmzA1uJLTBx2QiiAm/H3VSzMxcHTVy/KxUZKnDxwKoI46dW/AZU1+L//aw8swdPFHIrj0g
PtRo6fOVgHKW4EK/rkC46vLtkoq4jnNMaRMraB32AMWQXUU4Wy+wjTMS6XDiFFP/StlU1JP4UozK
fjrXuCFw8Jjr/q61oWiuqSM8kh7gcWh5Y0OMF12JKsuefC+Yt68pfqA+HWjSMoyEj39eUBpHtD10
P7sVwUCzHQTQ+yszU9hD8qJTVVhcqzHhmC4QtmLOl9WZvjw2hGzDThVWXD3DYFC0wJ4Y1i6IYxDu
lkm1CaQH9PGjMJuLgOsMRssLTDUp7UTV1q9vXoSB1U4El4aTuqz+uKUfFrhA21XGN6pzW0L3gr8s
xI9eJOMrVfuH6o+0ekih79hFLkn/7cLCv6bU4yV8nbG1p9U+5fpqNAFaWRlMrGeffqSMc/2b3+6q
akYido+NgM4gO/ZMtquL7t+RFrIJzv78zq5XAnN8yjW+jAKaYQnuGTExPnw8IZ3nr7fdKlYTwjPt
S7Zw8WpPwCZX//0U7Vx1QJlQpMbCcgE81W7VK2BZheynkCR043D1Na4QyTOtXz4HAjmDW3YeGfNj
9bWSaQ0SAeYnzNcd0wVBVQ0kvDCYlxtZBljcve/pnKAP/ukAGJRMoxghnNcwWVlKRraeKRiLCm7P
2hfaERpxBHi8AMID9Y6vGAjkhR9HlZ/iYpZzcjV9S38qnojNbMMpjEuni/uvjsCjXviF7KRYZVJH
ZUUs7259L1tJa+kWstGTaFKfj6rW+Sq8di/qwZyW9nFpJsUdG4eC9dlJRusS42zdyVW5Ks1iGWf7
FhoY1xB2JQiRZRwxqwkBmGLhsgpjFAczVbZOqgA14xuETBsdvnbrSVv6wf/ofRXKrMqFk0GFducO
PLd5N4NKWLGULVnlEIhSNrcXIAmPvON2KonhlMY0916OugDdI+Vyem2M1/P6oFILHPazS3I5fHih
8VEDt+ISanTKH3Gq/eyYRhhOTejx7Go4a7+/9pn5O3lyOkYhWBdFy9HMCm5AE+W5xIeYF3PqvOOa
TOCMn7w8YIa7WdzdweBRBA2p3YmO9PFPPCtHQWeGk0DMqyRRJ8D+HSBDOX6cuDsjH+Yk53Dsm/iX
J09uwBXAXRoQuQMd79xlKHHUDSmlLhSiCvQX+AsbsXdSbMo9knCcxOXeKcFBLwavcXyE8uxfTHfY
u7Zs2W2lz1qB4e42+znZcWM5bASQDZeCTrLolfwTGtXk4YOGBQCdVs6yxwmQFTZL9fhWyxgNue3A
FDIJRMQrDcVyqSug7h8zTSQ6J4QlULY/aZm8btLpmNgohRDZbL4vNZoCEo12ckHihqfH0eiTuq7q
jmmNaD9Eef7ZsHjOQqqW+7PASYYvyyzfjFbx7QX8cf9Al6ZOsMouKMonQqFaFHwCrlZL2hTlofOW
Kr/zTUDolC4NsUu+j3YURxxRAPwbYfwYuFjR5Q0lUlbjOxoauMnfLMB2J8kU6AgL1LYdEJ8FZSG/
oFiiSPVofPFndhiysw+p6/y/Z48ZUJAxKrUrQGmSimOqjs4gzmPOkzBTcaA4W/1CJl0Z708fYJRz
gp2JTP5SSZartswB/kJ+IKpUPLn7D0r5z30XhlJdytl1BbmKi9AuARwuTbFeoip8aXKJz/1QJXZA
gMVWIF1N/1Fv7JhF/5d1l6s8EwYK0X/9/wn8AERkEskjQBAoj0VxAFNUArGddHRrgVRvpwr4+aET
8QktCLs3c8eLPm45PlpfI4v5B2hGO4W41icNtmdB3E5/b03hWe1zqHKWJ3pARvI+yjPlXZoJEl0O
HmeZjAII5rJzOgPO9F27CUZEtQKAXuHYT0Flp9iYmgXhuCIVpQWBsP9rf4g88MwmJZq0zCuez1Yt
W2Ipzk392e7+SOXRJgzmHx7nvD6NlCRDN4oJHIYf6e6JgygGTkeAT/rg0GynThg3GBkLDZGRen8F
NU3V7VKMQYqtsmkEK8KACWj97S8sCmlASljX7V7LuDcrlrLXU96PD6X4iNoSGNcfC8dqVkg4bo5D
PpyEgdEvKEVvqRAEqRViQUax/lPbbHAOM1YuCQDVWYNCisrb0/TqG5rhMjG5UE4vU3V4CK02YP8H
Yem5EKgk1kS8kREXKz9ljlXMBmPmk9r9uqVk+4rB/EJ949PSgexpSlnZ7d+d4tV48evm4AM5DUCu
goG3saMq4V066AKFqFVq9L0w+gE+iOI+indK9q0M9/qo8p3TldU3yWUwWX97uRSN9By30lPesTLs
9rghSDl7PAG+MhcJhHLiVSZ3SNU2SMdMgELQ+jp5dYLclQMzEVfVnyiF2DGch+VB3UsoO7ql9QP7
XXWK7HjZttfzUG2IYKyeytH+B2ExKp4EqlShwaJ+XHd80cHlMLlh6MbXjU8WgvuSaGtVpXd2Qt5h
TT1Sn1FmfI9gD0Hh4ppDJokWpb6m1yWqoXbhmUoHX4fRcz21tyqaT7HBY/f7AlAw2gPknyWVyqhR
qyp0tIEDLI3aIa+zg0VuFu0IWwlusO5bG6jSUF3va+5LEgFzyQLeqmSFHDn/gA4fFkP6qBb2M8Wo
P+os1M75D9FC1qbL8HLdupsbKZVLXyq4mypkGpbyz348QC0Ej4zkULKVoce6i4L9RqpbsEEGILxR
iwrQ7fESoKk6UsQ2vJch580pLDw3Ylq+ZdVLcONfTVKYpimWc+xYMDO1cMyHKBuUSkZWmJxNKW+p
+ez6v1ftIUMZYH6O+9Y7VwadURVbZpczkEp3zjUtftCGXpEpIsIm/jhqqGp0ADdIhucaPV1eS7M/
4WGCXuc3w1+bsWeLYaZHWqzO8YKXDgcHDp3a3A/wrd8eQvCEDJeXDgB4Tpd7i+Eo6egfNYPfVb0f
dnGPq+8YZ8esz92+tQKV3fSnzuAFjrW+OVvOgIlUiRHExgk0dpQiG3osWa9g3GU81MnPPGg0K7vg
qJewd0Su20HlhSHEJbJamvVGipihn/Io+gYDPylYnDGbFgfkTNkRSRtax5/oAY2DYgMHH9FyJCGR
kCvh/xkuRc38DldgOm6VjG2VYFnUtB4QKxdJh8mAXioIrvCy+zq2nqH9Qh9WxRS7iJMzIMef3L8X
vSy2oQd9h2ePqSUGd9/BuZmBVFoS2BBOvYBkYh6WWgdVThWxonV1azUjX24f/CHI1H2TBuUPJQhv
tt4Bg0ZeCLPFC/g2JUqay5OYuQlqXVAfzvtZrMmJOzgHmYVA3lUcrfVOjIM4j/0O69iKbepbdTv2
ksdkPai4ii/ecuYT5cq8hVPFD40fvwfINRKAflQ9O0Nes3NbwOQ8voh5mnY2tcMsFZdDu1tsG/OU
vdUiAIvj7cCF49wgnFJ8NptUSVziOhDPjbfLH+88NnXxKiXjdkBZzIdKxFvNbsTuef2tT0ypsdhv
MPb+VOtdj2ZjQXR9CO/8KLu0w/cDzOVYu1J9gft/6QMiKxggECLN4Cqx9UbsjkrIlisZJYo2dX7T
P+stmSqmlPQcm8JjnJza8THIowKWpZnLON747ZTuyJv7RXCpFbc61tM/g8LZuV4030UMDUAzbcRS
CfO+NBkx6cuUwujTVeNNjtF1nSWjCcRCOuYNY3OBomRF+zi1RXwNtmL/XbFCYqXf7fYebkl5uPj2
yB2wPh4NuJyafH8Vwevp9ffqUHXGCo7bE1AFJ7Ckt+D0ECN+4kijswhZDZrw55CIJQIom5eiel5t
zG3lxI2JO3SYRmWE5cpNw6Ph/lT5QL9+Isnqvmpv+W0dzbSp+Y1SLX4sAYzbPov06aUlhwFs7PaJ
MIbb1sjAoBbZ7dZHlYLSRoKVOzzn1lAFcPMBkzOntkVFJ5a5kUT0ajJRs7DcNU88P7t7Ci55TUwm
JglEd+007CLi1VcDXERI/mIUESVfMqxq+Ym2qVSoIl6wyPwplrAs+3MFruG6oKGY7pSVDapodmaO
O4sNedCQnYXxGl/r5g371dtC3nLOtqM/RSD5iwx6OhDuhnal4iJVa4CfH2Dq2ozWupiL7eGMfL0v
V91SD6fi5Vx14ZkIFe6u9XUR7qsmXQ9TeNxDFGnAnNDT0aTidbVhqpxnv8+uawhhIhTXz+jBOzzn
5xJiTCD/6uO8xuypLvXykS5oR/Ltor19rPxqons/tMXi6o4FxXFYMbhlleMfTFoWM/zUc0Lsr6Ai
0o5q3mnbhPwxkndlDDWCspAtOfnxfVAg4hhxMzTX7Z9EFDXDa08gWi7DlnOs6QkGeUKVGfKYopn7
5QKUvFVoY/xjnZQF7m49yGq4BXYyZkI63neXsINL0GIewuizoQ04Von7J6zpGeUwk7a0ft/IH/m9
P+9FMT77PgliTogsiwwRK1clE4Ky9TLe70IZs2ESW5EOGOEUN02tz9ibe7FiMS64WuLfGhMVbgMO
zINjwU/2ldyQpsSK7mDupnY9NIiHNp8Wep842b//MoOVelGfnnTT4dB8Ytj8Kq5nB5V7nEGNLaMY
bkUlHWGhWlqsNJoz1LjMbcDFNmjJ5fZESbg+hjeTD2dVmS8TFKTSQ6g04o0mleoiPhO6d1Z+LpjC
mwzNUU8FSFC7V4wJYZJgxm+1op8JRLeNDXLLh/vRrHn5CNvBCUS45cAvKdGW0i9VHGYaatViUMrF
6EX63S/Li/Mp82K+UnjWlvAZCYOVIpubF8cdoeLlAuEdsQhSI434+QTABfxqIAPRJv9T6rTf57gl
7sOpQMtzG8Y7PoagjK2/1CIVvKeJ6f2nxH+BFeQRH7KaE+EpGKjBl584CAm4KUEm4/eYbVIV/Y4i
J4y2kvFj07U5BfZ3t0YwSBtC3fqJ+g5NaXH1Vr2RkoQPBRvjPiD7zb4DyvUtXikGDTJLNxRtiQn5
e4VAaNOc9w87WW31vZhuvigocTjqUJj2YFTggFF3is9Dn4XhUJAUk9S0AONtjpW0oUoOEPPkRBEf
9DS2zyNPPqLA7CHt64NKDQUgFzV4HpHOogmcZX0KB8ZEp1RykjZGaCk3UQA2m/LI8cfajtvOhD5T
wbSZxvqdyvx+6zTnITqLdyDGqxLnRvWEPTuq5u4Qq5aMnsAW7XLdzMapHHIU1uGwf0MnisecZlya
3C5GfPSQ4wE5V9JvegOVdK3IzdQUuxXtXjwy2T3xA71UlsYBi8OlQFhmGhzjFyejn7FjzoWCR6fY
gilaRxwC8tZcPZYdCHGT5Tf/nXtjDn/vXlzErCoxXdIXN29k18QySerVcg1pcHQ27KZ166j9LYRM
V5k6tH4Uf1FznVyDuDnZYZSt5ZcV/O9+YQ0BTF1R7cM5SWCbC/Eh98h6J0b6bg0cOds6XacBu6b1
TsjXHINo0Tdv3foowdE7HjT+/qhGrbgP+7tCMj6SRFFWQ6Cho8Am5stiMEk5PfoXbLSxaDrEUxf3
xOtoYp84ZFaWsoHC6JywgJXhdTJbfJJ6drCFXLQqXX45wvqiBM+ezPx+lg98WJAA0divnd/qOrlo
Cwz7hO1vEB/E7wXVl/vxtW4qWzP2EVyzWzd39wzevLgHMo0AgZYqCokiJin5T7Fl4UeRa8ze1NGj
AqBCHMNkVKNnC44ePYD3M80AaCaxvgETUxFtXuHXfK4SM2QNpt1vpBPfBarUjsYaKXDcTGusQP4X
168CShRzGj+6G2LWVtWqzdS91o5+op36OCOZjhTFZN3uI5PqnykEmEDRRKd01D7TLUGA7zBEFMh6
/GmhLcKcAYGmPYJVF7Sne1QQL9zv+OnsnheMJFjQX+rTIPh/gHlERPdPNWAaPpwGvu2BpAyBE+QE
/sAm/7altF8GG0xDCJeV1+Jq+/zwIZjYElgkP6qU9ktEsGggZrW5GdVo/uhNBUpZvKrlEPWVuzub
CzjyplFt/YFXbMEga6KpCGrNoKmup7n4CVKNzxgONEH/s0z/wvCGcVwkv59Hl8n2pkdwwtEUFGcM
xeJKX+a70oCC3a1p7NYkg8f/wCyWCs7kYXIlhfqFfpmlRtjk8e3xMmVZWk/I8R4G9SkpbPPDxhT1
Yl8p5fK8FTnw2OijJNAhIIE0iDNCEtjFH3Inzp1onbgkehFzfh+Wskk+p4pL3w1ohlOAfvjOswUH
3/ZfjGSwSUU4tuk4/EfDytjKQMbDm0pAWwj+XlOYDZxM+FX+0hBLyhuHhTGHJkDcbOaia3pBUOvS
iWqPbCJA8x5CpHHykbaWmKTi1ego8F57UDFohhA1D3fYc8JP+AXAmpigoLG+mNgxCk4aNxGyLFUT
P2mWtt1/vkhvnwPM5UFYSZ/KgyTRUaZzSA5CbiyDOWaCefiKNcypj6/jmQWpEvPYICWHBpsqrgSj
bqfKEit9IJKhjxQITQixzUTealceCrwxLSN8vYKe3Uthcv6KlHuvoQz59Ro06ALf0zRSiuy5yvbf
6u0OPAD9rsT/fxtPHRsR05O9UbY7wIz4BsQNq822P+81KyuGNCHTz60qOPahrs/57K7MyD+SPMCu
hp3fdnbtBwKiA9a8InKBB1WIwttFA95kXZi1Ugx2457kZ2rHwMofwoc89mX8ygt7m0hd77uZWQPr
EK+khtFYOEDiBD7s43XKol7N+nRIPhPYgiWkm+jYr85e42m2ef5f/yu63gbWBInsjXyAMiZb39TC
9cm23SA72C3HkKs/hfHZ5ljRZZyqloinz+EbtOwLyFSENuXKjvkXsXcuaMuycel47egEgXUhq6mp
DA758NxKDVNipeebQmjsadoP5F9MwaZfhUwqXE3QgX0KAbsqsC+OhPa/Lwo9xjhwZChZ5O9vjFTd
Z1i2UC3SZWn6FVJX7W41pueAzCvRsCtXTgRxIXmJ4u1AZRaZ+gCLbBMmVhX2mMONanF0PO1BLJMr
YsXIcwF1PKnoZrCi/5ox2AruVYcMpogt/kccM+2XqWGVWDIUv//UQ/jUOWVWO/mUlVdFrlfvuqVL
nveDeRMuNqPGzXEhoOMwKt1/88Dmrhk2k0nIJ5hyYTG7HKvp3e9SHQrZ/y0lcFB5q2EsAMM1LCxc
T3WMx2kYB6wzHRSf/Uhy2FLVNqOy1pWTH2HcBJfJcmWvM8EFL3Je/PKV+1mFrooRJkAQGGBuSTr/
fsUEu+YeJ4wtD+kkQSigC/wSrfs7FhO8aBWMqZinM3x5bXuWtmZXJ7bIRuLz094P3WFnQ2f6fBJr
ThW4xabUk9lWDM2Ko5RZod3p5o5o59ePMS6i9y9og4bQcsVAuVjrmy5n2qBl7ioH8FMB3YLexEzT
joAosv44NP/KsNwsrv0SenTLD8KmzeP+hO88CUTm1lf0iFNirTUxTRUn03ol16nZCvGi8sKZ6vZT
z4WEDIWc0R2iWIniZI2ev9zy6h0ZwPf6xUiBTJLf57ABt1oA3dsSSkKcrt+eLuyOn5ZcJiplZkPx
AmfloZEQO2Fqixm+DhveS5Hw73bV14eQsw+K6j/cKQsMM4hMbuL0IiFrR12MXgaxqiZSgzhKm/LC
7T64KTkIRVp3873rLtMU2dQkIKpxa3fTu91uE/RrV2alnaMEbEUCZwyjeJ2QsxgZIRcxQDKHwh5I
q+kUoFaEXqkGVlxlSOyD2RF4jihKm+neFvV/VI+qnhx6cIgfGtaFDxJmAQLUCiBJUcmmIXe56o5A
JGE6xqmsHON4G2GZ2YD3h2UUUyfktsQmfMcVMmWrtogpdyAj7HTwE2jtdMWEgannd1qT0Qmrxy8r
CLXWteSvJyR2psfe7zLxo4U1c2kx6y0+GEk9ZNj4abbhehXXJ2v1jZi+MyZYoAwiHKMVUuMtEVcw
anHj/vywmFuvKONgrUnlXxqjo/l+EbMi0I+tUo0/h0wP6+1Ncb8sE+Jum/v3G/yDKLWFF6cPo/L9
3hO+O0uL7oPsw/bT1VGTt3d1bskZnQECR21sTbWt9LGHtuwFpFu1gvEUGASv8BYQysrJmD2IGCrQ
r9z9D4cx9Coy0eRZBJ1aVRs4q8gWEA4SroBgQ2rwXklZ309KbcU+xoF2q1q9c5cJUbxN4wQslFCi
m3P8pXtpP47Q8PcLANmVjcfxs4w+Isb95M4IwXaOXXqHJouxLJGCmesxdhEOYc86McXNHfyHkuoZ
EroCxcu8+KVofLT4JFd1x3+vxktc0q0racB11rIVuqJrRs8Fp0CDtqSuXxrxy2Zb0pfqUrMKto47
sEWxGyshlm8bttWpHRa25SeuIwODIWIYc9rQTkXq57CBHWzKDJUTbhwZ1LHjX22JUPvA6c5KEwxi
reprnNOlcUmplntMsvTO1zo+sVzNgnBOnkjB/VTy9nKE6KAsa98LxNZxa7hOn+4qaKPjY4nubba+
QlsNJbXlPinDwDZ9+evmnadn9qi8MU6BjAMtOk+pwCmBx5TWtUz6z1C4GPO70kDSpgSlKsjVCdG6
GYsrorqFv/95Pk3jLEbjZsYZ6qlaRoLvV6j/dziYrjOXpI1MdN4Po8cW2Q2my8OixqY42VF2LZ7x
KRz7KY8d9VpXpKQEZDntU5xdPSeEsTXi3Ov5Oc1tiLjDXzNxl050fBE1gbZ/cbGhQ5H6b6p8eqZm
zJyWOD6sV7z/bX8CjHr2I7waa4fuKKxd8UqVLwo71AefHo9n7sdxG+RQqlCWSZjG2V1mcd8vdp5B
D8B5sSvpYhXZ17Or4Qh4a6Wg/pPUQO/VHHYtTraMXRlheYXC/+F12ajxFHADMPyIVzNQ8AvjYvvl
koNNBzb287+MF7j5DKWhjHod89/BByiIcxvXJrLtXnSIodT2oTpBy05J3UM384rsrbmhwXMKF1ky
s/whMEzVYRq0j5PQfqc2I2riTNUebC6vwVoZYs33Q6BCPwhgMigzx0PitVjBjOc5VFQN9JQVqXg5
stv3EvsURmb90rVN5M9BPyOoY5nySTwSlkzW850SObEm9UnWbucvkaHVCqPMN1w/CjZi/+ZF59vd
oIUviT1ak2T4WNMBJxloGvMNhNSkh0YmTg1vUS5tsX7sijYpuHlUiuicwOGrqew3TuviHjRO9awz
B2/GFIGA0tIk+fHNcy2/Yg9+mG0SFSte+okP8Q9g74rxJPmdvi6pnngFlJQGTpPZvFRvWgIFglQr
EEgCpOAj5DJmE8FKxWwazbp48jn9CmVJEUdOKNnnI6UvVO/YfOKKx2QSCVX0Y/nHVEHIIlNYK1Qp
evSQ8fHvdKZu3TA2Y9Qx04IDJfTqRomChK3NaanVKyI8KHYLdQ5AxAVHrd0caauK0ZfgoTE/3DAT
6ezEMltXfDJZ4jfHps5HcyDEgGUCyfWJpI7fzzzcLxEROnly08gFlK+ZCSd+oX1XMTljYzlhtWdg
40TOpk22RfZBQ6IBsu8Pqsh4gDVMXFfFCCS85EoMLUgPSLOuUU+sgwPfmgPOAMtUMvqRAeaRq8ST
xJsOudIGnDcWQssVDRe7A85zkiGtXdogTd0SWomzQWvyVyDbl8cErCk0xGA6kw4Qpb21wCL0dWXM
nhzmBLYUlPE8xf97TQC0eNamzy2ZQnARp9SETeD0QXbFk1sEcjPPbV5aCex7gN5Sgy86EVl85yuZ
JpoxoBcVLEHPpj0xN8qeZ22xDWXSxTjnaEHwN93z2JMhWiDY8EmN/s8N2pExeMAIDQRlqyA5fi2/
82OlQKlmwuLQNZFSZEPEwI3Imhzsx4RviplmpRK0quVRBfFnRbONMmd+8jVpd9o501fM77I+Z1gL
6xuWCf2oM6k2JLEnO+HcOJJSTZ9J9qzQUuMMEftotCswQ9FxUIm44wK4ZtuV2s7AObAMkFHSd7Mw
NPXShZfgldguXXaM6an2FqaZJzhcZkj41wCCpq0rWCFyJgGKC8ejyznVLgtXqdWKOYAViUEGUCMt
rgu4u3itV94YF62ek008peb/1FEqkimv91xCCtZbZhjc213Jkllfr0Kr8c8qzhAotUhoEAS0AEZe
G818zlDO0AHrGuYbX/kvi60ICmDaAYFMxksDKq6ToBImE4tXyQhAUVzmmDaZlgnAabLz7Tox3g1m
LawPfbK9p/C3Rs5bPOK5guW+DdBSyqrfsw+gdjL6A0yH8unpR4tamdbnhoq5WAeS68QxE2R3iyg2
PQo1LkdubAtOhqUx8YJQ1yHfJGsN/yuEerSV8NlRE1mUDSkB+LEmPkeH97fse/O2arqKhQB/xyPs
Vlssc6nvs5g1CZvuGP3MMTFuatgSZwLJ2p+TB0X6OLDpfgIaNLLFAEwRoNPuhGyQc7fHq2lkJcrV
x8eT0OTwJnv3ZcEjP3AfTgepsG/DjK9XCCEZGO+cNdY6eDAyA8QH3OxjRBHjphSgFtsnmnhI/eC0
r6Dnb08Ema4uKbeDKrH2Ct7/Zho71PfIdyZ7sG3tkSlfCqxROnPCtG88vJa1/g79qAqT4IJCbQ3Z
/wUa44i/4eU1HKwF4Fb5CkS6A20Axh8+CWK7u3RtyaCirTR5cOwTqiEUhQUuapTuE8yJ90b47fsC
ALy0aC0Z2LbKzvNTmUsMFXAA17w/N+W9vTUnHcdfPRdIN57ULUJ+YT5phx3w/9wG8IRVBkV3MJ6D
TGar9GkoeOs5WbGrgctr+gUhSEz2HTN0xjnJ+Z0pP3uIgN5s+BcylmEGEHezD3eMOTgiatCMqvGQ
I/f0Bx4yRHh4WJgsA5Z7a2epCRKmju/UiHPaadD3TeZDeeBpSoKWH5u2q0m0pzoMB4vA/GDQjPtz
pJWMHMnaOjSDhi6hk8f/VcqXoqNz5L0/UcPJx8GcZI0KMpGXEqnhYPsOQEssKpfYxLUAleFvBS6J
77dkTQkV+ZX/EBrn8HyessG+Wv7fxGNPNYWzBNX46tzQgS6afg3bWLlAxuDRu0ji3eJ+uxuMoNfr
UiJKupSSTR5+8fhgyVwlwqeQu4xBzhvKDVvJIEyIR6IUjxoyqRO8iVudhSk7uoShvsC+/ZkPGLKh
Y3rHJj1gTwFkhkFYQHWVAvUQWmPC+aF25BLuRrBxFFdUgTKXzYSpPuR7Do3/kAK/tWCVpM+tDhY7
NlmRQWY56dMR/OlVwD4N3e3aUSkp4wogKcXH5SdPRrGJAtGSffetEd/CGewHqJSqz9cvnJn/OuJJ
KPhDZeiZNcgqDrdbAfjNMOnQqbf7vuRPqbPPcoGkXpdtzimFJ4aUZDA+zULeOrYQdPsmiyYzaz8P
tJ7LQu14pZYDLU3nzDgOROmC7ij4tyEEI23fM3LKSZHDLR7s5+Wr5QDb82ejI4wB6j753inR0LCh
yGggqeVnJLF/+CYiIffbd8ltCNc0uBmjfuiu69pN2gkO2R1De8k54l8HamIhyPDdhd4MyjxLE18z
+sKayAljxLQyIww2nv/vjCMp99illnDsK0C12TYP/Tsnw4d6kQ8a8Z4R8LYMg/lu4Qhf84mxrS1N
GUU4E2ITkLRMvuTWw9emqfcLfSY71FhSmyG7dCU7Aeh4ggvgl47xKikdX6uMSvftsalWsTkWDiS2
IbjcbABvPU8OeE57uFecmZ6A4gUyChs4HzDkqIceOUECPssLcH45gPMOyiIKP2H0HGtIUj/C7W9f
iRaLOoQ8qTauw/rPlp7075iG4q8VRSJjnrVmH2VKNOjQO3Zyxk+2UEALjclC0PoYHas414HjLoSf
hLWe9Zb+yghyXdaWv4/vmVaqtG0gvwDdnNaUFUleTbm8+NIMDOs6qy3amlGX5EYKVg/AhbrDNV7Z
VLPNa4OykLkATgEbBiktp8wJsQLTgb34gGKyh68zCKE50xtQXrmDxOb4OUhifwAb0ZnKyPO6ZIYu
n0dWF2nkLRC2T0glfU8NHSM9/u5tguP3cIMNE+4EDg6Yf/+6+WcqDAMNdD10UUhBZJnUq8tAYRZs
fEBngIoX0k3C30wpoy9SqN9pgxPX31rDLAO6xuRGhYybXgD8Dt2VSNbSCAWmuWzoxJU2r6dM/hPP
1UmS4UwEQ9K+rlXA/BFGl+Dn2jI9Ag2Usue3ElGdavwSYlkrupNFo8b7O9dzcdm42qNHElj/Wtf/
hMRBtcLz1RdjB+czuLl1eADAhnzquI2U9kfuUVWJmSnCnI9rzIkFGN8M5Hgw71nSpDfMiiEea/mv
m3QMxUAz9Tw5WeLgotcALbiZH+RL8QXgvmHxtt4NpFD3Azikr+QFDIQdI9mo52t/c8IgyCM4cp+L
KXJsdeODCXRMdxRy/i3V3udrFKLk/132F/fWjvAneXbnwCX6uw259OejUgyBsVdfR3dVodvbqf1R
Lu1N+XjrGC436VIW91Abm5Atv3K/yITzPwB2gXKJ2wsWyR3JEIVko1cpYVLlTWUc2NDSV6lwbry1
5rG/pAwQQZLg6Y3e8Oc/re/HXwggwFhK2IxSVcDXJymidYVBorRp1bMbOP/k1sFjYL2xHoEr5J0O
ddGgKodZmKA/NFNnnyIqixlHiKifycfQ3ks+HFP6KU/hM3n+85G8TVuGsHOTSTPitTMsnkf1zVF/
y5koBt+Ti3P9yz7se4K3wXW4SQS1ZKcb8wTWUrUeO2NcY2H6L49nDr9WKqbW1TLQ3LyQ3gIk+0uM
WUh5k6v/l24gOcIHbE04zsaioeTtLn3rPx3L/4iiyGHmr3fq3zj0rnFTgAg6sTMuJK6I440iRMmr
2kloz6BYbT+DXiXpIx3v//ndHcpmvu/vCxwtIOEm1bbQNNUtYJQ7ZoFpqDgqVgxcJoLIVv02I/A2
y6ihHan6vMa3SaO9yocWGnUakMUdVu+n1qqZA3QA0IxZS18FTvBFjz5r2h/l8MLWG5Zeqrn3wpuE
ubDAYStx4nwwivmJjlqevtd4Q3H+Sff1f8e9fq2WhJjesZxlAqj6K/zq/iUV/e9oHBeVWMjVCbLG
B+kh6sZv4AL3zkJ/k50hboCgVBZ10xzbxAMLNZiqtLTsdVnx0MoPpn7uHFeGr+FLzF1Mt8Ggi+Ls
xr/WlzlsDtekvTRhtrWEnkmE1HraD7yrs1ooH3jZZ/L3mPMrEVE0AFlcc48SgucqGA2mONWsSDxp
NUC1Vn48t7CG0AzBP9eK0Jad4lucCWqO1nT1O8+NpRShMigBGsyl1VCN369WdrNxUJ+kJRpMvnPk
mXoxqZEpXxDoQ8kVoW+mJYgFYXXVW9CeUFOeatgsSB44gjtlenY+dgjSu+8Ijno/LgzCVJNEs4Sj
dlo0zRX9j7pkrTlSwg4ZmiDvYhmHLxyYIehn9XPq5J+uo5FNx4QLUg48p1R+pgQnGBh+9h0q0+1J
eRcFHn7CbK1RErPXFCtiwy10tQURUb8mONIRgwbwhFCqh936EPS7UladsIOsVen85qGFbCJ+xe1s
f7eCQxDcx7OXdNm5etsAsdl03u7ry2PwFDTPSZNy8dyarpVYQzq8ObZcAH5MH5Vy9S0FMLIr+qMX
GBDVOQFmRH5fFBR25cDXanNm72SUqozBUFUI+8NrJtWi5ey41cJKY9Svgzeh3dTbG8F7hcSWTTsh
oNQpF4R1lRBGkC6v7P2QiNAgyN5eyCrfnOxeGRKesWoIc+iSDRVAPMjiPXHUKTTnpjDEIsk3WAza
bDHch4HK/685U8rbHEOYzQhOX+04YfyBZxyDruQO3oWCRWdBXf7/sDSU8WfUn7d4gfI3VoAChk1x
9tI8wLmGb+2JFBPT1x0f7QlxZ5Ts1jTPcFTkxgwqyU/i11iM4LIxTJ4Knkxd3LrP9lAAYF9+ZSXw
1uy/tUGcTN9b9DmVwR5CRG7nrMjP30SFmbdoxkSzVcZtrdJfxcPSFxSxwXlKV6yquWFos5iePf3G
Ue7NlPzv3FOFOdzyAt4SPM5uSbPPEaGYoYX5BPRpffUDim7ErX4uc+2Mb8ok2r3l01FHF1+KDNg+
K8pJ9sdisKqrHvM4rqkKEIOuMLuSVZeSXSlbIgyY8TrDyZv5Ltwsnn4itxHB0BB6/A7UGPbTMZfu
7Dk6eqUiy7FwRDR7/E/uwwdztkLBgcMnuNRD69e9cyPcPfxjruj8SfVglyFkmJ5hq3/i8lKGzzIF
WdNd/W3l4d5VG62uQcH7ZMCwGHoK9RMLiAKG1yb2TKo7gK0qHXO4o1HkIVnVRlykuhmjG2C9xMEY
YU400cwAwtwIpmBCFBTT+qyIN8KAjnKqCSDOl1TK4cQb/0iKJkAtCRUwErLg5QhDPGjzZqvqx/VX
tztdBLyx8/1BKQoZKrS//KBJ7fKoVsdtkH1wnG0JlnY3eXMZ573YC0ED3tgMhRkyckG6kIUE9Qt6
1pK2QIQwg6JavBC2HTFQsUn3jwQXgvhoQ2ma9j89Ums9VWI0xxSKlM7N5BCYCRd2R5rrFHf0KYXL
UV8ZNTH9BMuh9qXHLcJJFUZzqnaYKS3o922jfPpCoyaX0AiE0vy2J8AzFU+0UG8DAwvtGNdlm8tj
qMs2gFLaVQ6FlLvShOt1JSzVANE9PYJo2IVblm3eYy/FsE0YBtn0zmnVSpes186ANtm2ZQy6imNs
3UlqDpqReDSyYhsVjLdKgk0GZF5tEigdiLRaHxvYgQj7tz+0sqYh/OowKkTaGqYSXyQCCS+EL6na
WjIFDSfam+q9HQdsE5jha+DmBwRlw0C5G+bpMAzp76POvn3dxhr7vD+hk4xnFUdFe9oIow7w2R+T
nZLbBHQEyxAI1EDPd6ngG8t7XsY70JymGKfvreuhwOERIpDQYPbW9RL5FeJ5B6m+pdrMx6ZGFsCJ
0bi+t+cdxw582HkcZNHyi/bRddcCLUgHFIGLrH08G46XQCdlZQEDN0kQbl3N36YYsUPZizqZcRTc
gLJc1/k9xVGB9RGfVJ+yAYjs+d2u/hNZT2h8b0lijO8X1Fq+xw21woXMBNat4MZuIFcNnHlwx5lu
JOU/K5t4pcIqD8TFa//6OWKWec8Pidh7RJNpk9AXvVhVqdfE8UQ06IspN7fWZlIDsksUSrXcQvon
T6G3oz/WFv6pJwabzNoAg7kHXC3tDDgEjkw+pwvjZqlvVyvP6zl/fTkMNjSEomRtAn/07l7qiGHc
tRTdcarqF655dc36C9WTxgubZ1bY6JRtVj4R4nqO2HdmFCSd9IK2wxaDQJuMrZHLnrbM1Y5pI2yt
a+p7cb2BLZGp200hc2V2VhVGXZS1OV73eEkXW+0HW9bjzmR3C+19jRKZJ1WNaCOeUPSQ5rmc8yPg
wdi+jYfJRw1B2Bqd08kxAFosnzmV3/JUKH9niPhdjLXZxswjHZsFk5OnesUTOwaWrIq/NDW7yoXQ
C5KMLNyius8440NZzvtvH/J9m/2n6hBzGy3R+1issgkehxfB/efXwR19Di8P7cFxO/TSu4hOC9Iu
hZzWbsoCpDonF9yJxTshDo5LZkm/XsskS2ILRpoCZqRKguVckGMN+ufF193kZUH2PJtQDiRPUTKd
GwzgGqHq0Wur/mbmjir4EhUuequbf8MVxt+GK5r78bShh9f5/CmtCqbjdRC12r+meG52sv2QJm4v
YMJMIYAICQNPalWso17hYjq8EZtZuL/abh7ku3fXHZk7tFXJku4epzjPzIaRQcCDX5YukjVZ6ljX
UQZeAjvN4JFyzDxeKgcSfTPp70eaqNBVt0LobyoBiWa8rBD/upErnc0fBQGsnbCOkBUe4MbfpL1W
RBHG+p2yrO5HbIS2zN4tEpXBwCsqLf42kDAx1+DbYFaYVX1xIHymjwmhMCGILLueMIccVgZIfj68
xUCmNt+M/OdtdL/uFBfSwq6/2CIHQHcOiwf2UMRDYeaG5nOY/IkPQ9zPKWBRkEViVVBAANJufu5V
kYiZO3LaMFrGYaY/u4HiZRs7AuzS8WoD1NVF+GIvRmLVXh2shUArfLcI9tVN/NUagv6jEfhaSLKD
L0Pzz6hzChx8Xk2AZFSta48gqXgDhDrECbM0/4nnziC0ClQACKgE7MVKTsdDGtVd+O5k/bX5NrJd
nXLMPP8KrrpdbYSbRE6xKQN/bP27obwtvH73V8V/7OvSobKmwoHq7Vbk4PS//a7Ij3CMriSQ/cGW
DrW1nprv3XRZDK8iuVbWkUt37B/5V6VoeMrpYLTncwEKKP5dqxQRZQCt2QV4OuqvtbxxDXyEPYEF
rZ99FdinQuZs88c12p0HQd7/oG9trcy8rtqXB3DfOqLaTQkoED2O1h70ZFFhXRYvLtldNzgD1Gb4
tc6oQzcIyn596qd0GUulnG2w6HQ7fTU66ir7ixMTd6+VtT2L0JqNZRVCSXSbgASkfCE3Au3J0H2i
mIAnrg4qIWEpPT/omnRAlgrO+9Y3ETrCiN+zgxNtv/bmmE1bfskdveRrb4YHkQotV+/iqb/KfZvA
389DassRaWn7URW4PfxgFTYRKGHWhzR08bQdTIq1ZqZAHS0Z1XgStD7NdPOJGmD3YQPwXYLA+jsJ
7zEgbrTAM2/SbSBp0X9MLRnmfnjY7+oMqGVMExPmZ3WeBXfODW+5HlRST0awq8uYWbbCvlGRO0MA
ziyxg6/FLitCVWBI2E1gFr8kgoJn/OEIvKBtukEbaLchxqToQYQ9vJZwcaRxI9Rs6mYqDc2DRqal
SZfnnWi21Q+nxCQ3oozvmMBiV9D9PfJtbw7YW0VgLKzAOt9HHkxtQm158dTgINyEuZGnH0boXFR+
D7FVBcyKxcPW9211WxL+QqUAkRP9ZXfCQUf7GoicjN5+j9WgPydIo+YXmrbUdVjUKGO9YPPFqOuZ
/i/uBjDUiM5OAf17aaCxiurqsvG5HhAPaFoHRH/r+rR4lMHfEb84mHo8XiodTr1+6HAhdREPZS8d
D0XhCQPlSK4wfGANDB9ihx9Xundm60TYpHve6oJT+XR8wzuK1y7VT1/kXHLBrOMu3gSuC5mr5/kR
XdeUtbk6epl3vK3GtgvKzNstfotNy84MBkpJ0UmW0O2y8DNpbgCCDCMO0xLNz3KQNaIpKoPtTCEa
O3TKpU4um2iDII6Odz3OHJr95WVTpqumf1aq8AhWgkTNOhlnJWJ7F/O4L/9se9fEJbEFxnF9mi0B
R9VNF71sPG7CnOh4pjuWrgClL5Dkdc8YgXIBy1c/kLqAYlVvExF9Qdg/1C1yHhTc2N/wOgrebVnJ
ZI7VO8Fp5XTfP+h5jB7GkA5hfWEzCsn6yuk+g0YHGwWF6QdiC0sHpjq1cihKTKWCkAzIA8Mr6zum
GYgYBFE7uCDkhaKnFiz6ZdRXHsxK2TeUgCnBdg+LFpNm/LwrHt8VDLuyoS1+da84axuo5upDaPSZ
fWH5ypPuSpgEyHwytHhfScZvISDkr8Ew02Q+vDUyHQz3kkyxbzoIoFYlYUulMeBFEWRjEncQnA4k
oI/FvQzxmlOGsV9VIH6u84U0Z4bqtz2eRenxFbmpKeaslgFcDWLShEwDM+WIaOHag3vDPEHbpCaX
SIZwhZcHXU3JgkzTlyewLJ9Zt/d/wiO2jMJhRNPh8itXYzg4rQqCSaVfhS3das4JL+1RTy9KkPxg
7+WQBuOohlHPWiTkkfe7WI+xVV35mpLI3j0YihbIeF498cjC4jHJj8USpku+kUddIGJPuzA2Vg5c
UDa0Oqk1fLpdyRcC5fW2R2OBDfEZlcltjQ+1zJ7LulRCS7ShRFxegb8UloZxY0pOASpCaF+nlwk4
qrORu08bpPsjgYJgBnQPYhRFWKzwbENtu3DnDniFgpaerRTmy1Glf/9zNpNQhxUPawZzvgIed2IF
jO8mOsuO39yIB5p+Arf2I7XIQ0JqJTsM4dbdNr1xdJr/eNscyBAfGLuwZHLyy3QzUy/uoco6ancf
L9tGljIcy8pONLTHuDeGMSHQ9K8mcwAmSSAh+s4Ay1IrKkUmfhjLMYRM2O2GlJfHN3QGU/OjPn1l
eOqxoxYd2HBUA1XZDRiFz/L+h76VsOAxFVzRXWkwerpA5URWxKI9GbTFJ0WHuAllSH4Fqa0eGqJ2
M07BoGUa0nEAXCCj0ZA/tGncZeAR0+VUckot/R/qS2iol9eMK2pUXd6mYNR9CKSIzu4V7LdjK2aR
2wYBoI4+t4XeEbFE7IJLnV3+u3BiTuqRcclBv5MRgSl9edW8nO2ypqEjaulC/aJtEP50rdq2M0bX
CluJDviRgR+cWIfWloLKeHSh06EXPsGUyo4pQeM1NZGzmBQxhrjPc09C2dGl0DKL7PQyA+HI3ffr
OzxKNvdI/FBHCBjSf7PBUouhp5K7BKaKGL8d1Yf+bGeFguF1QzfbLyKlqoSUbX7t4wuqfvGa8ZuU
XWAlFXIfl9p8uy0Sizsl/ti6b1+Csiy/EC7GhBZEZqQRF13fgpHvhVpVLOxR1WCq0ytNwm9jyzre
5XdL1gUnfcDvQP3SxzvOuvqzM9OAebP8ZaGd33zoxag2unHpdmcJeqtOp94PJzxhTrU8VyM6OZO+
98dpTXVXkl4oKUuwAzAzM2PLwTEgox4T/43tCquVv2fX2AP0yJ4lRp1dbpCq0HwajuqGLPT/8+mY
ad5Ko+rVOf4zAtIngbJ050GBV06s+D2YfdSCdPxXFU+Aw5XedFLZLjKGGAZJeyLbJXvJmUYQkWb0
t5rMDP+NGNobeJ3oYXLA1ECFWoA6eD4SnI8c2ehrnPUJAqW18h86aTcOwzu03NiY/WzdQRJ/clc9
EfxOb8BdKbj10KbFrbvU9m/LME+S/R0qUGfWL5c6CqYAdYLjT487JMikQpDLacJPTLA3Tjejya7P
Sh7Dhu3Di6KgCKFkwB/u+dd+Fhx5jW9KWwvHOZgty5bhpfm7pZAq1JCMMeYrmZEk0+0Xn2A38SCo
a7z7ixjMVJ9CKx/HXOgOoEWGQ2epOn9B8n3O7UFf5iNGZWNZIobIbEGRKoDPF/6hqWLzT1bXpkJ9
nJMNWWih+6DZ9tKUt9djqe1vuoypqV3sZ5pPzdNzadNgl/p6heHT7NtWOCTSiRFU+3ZiGrKGdNAT
NZvAmmjHXEtwBObWfDhoo7HMGPHQW3qj/iIzIpackq3bfcqoLfhte8QY46AlgHLucm1s8eAP/uu5
aOl38qQGRehcROBsjL93kAhmRNxvySi7cyrN4p7K9Rej7AHhpeV7JRyXS4IqliHb8Y8vGr+QjkwK
MGC/mClpVkoy0IimWwzSjvi4E8h485EPqnDBIYOCjb0RwJ6IIiOWczHyZIOPhizAB42Zd5Qpyne2
fEjUKvpwIKrmbPrKpIAhfalWrRcw3h7+St4fjMw25LDskfRDvuc0Z/wqR5adVNRiBrnhON+k9281
iVIEb0s02Een6zqZVLegugP1xE5KoSUsGbEDoImTa4epb4SCAIFLAgh60ebNaCFHoRGe7LQGOCoB
MBcuILmOZyWcQoin/zXmwNqAV5CGZU61FD0OIscZiPbSAOjuYp8cpxGgIIG9eULA3citS2Lw2XS8
8qaqERQwP0Sj50UgnUHuh1DXqrmxNxkmPW/6fOZ8cfBiUyW836EL+bomBQxr8Te80BG9lqt/ftBv
KuEdTD1xuRNwZV/r6rrH4flYq5+rdxqvCTewAN02Wp1F7kECl4gQMt824jo5jkRQxLXyPQRZ+bQl
5I1vhw5Zdq0UVybqSKN7CevkSm0Qxg4HxTmmQobMVxlPZVgA2MdQR99VWz4ZExfTYAXoEXuzVRp2
KG5qSaTchENv1wrItwNLSYqla9XXg99Xzfok0YYnGGnNlSeNW+8Q57Ww4ZRVPlFRh36smHwLROWG
7YBafA3ZdrN4RyliXnVQP2GX1wEM8VtGLH/LMMenNwdZzXCovDHqZ4LU1sNa0E3Lg7QD6nLb4Yft
fd/dfR9MzVy0Ra7zPKkUIYxqPC2tNuEUxQGGKaU0IJbW5yaMLbERjwJg0ZNd9UXh+03wMhzGEOyQ
bcNAYJun0q5UpRhlh7Ml8pNMa9pblGn1GWuP9EK9C2R7RQHenPLlBr3r5vApmqnYL6QAzYTdQx6g
cnTi884yTJ2wVoEwrjrnz9kEK9Oe9K1d1+ck4y8Q4hhXOtGbTa1u+93GAjWpVrjZHA/FA7oe5kbA
XyVjd+/nuJw+PrLJI1E4l50tWi8s7KSAXh6nhykpEk8ly8BpBDbH90DSBfQYDIherRf+yhaNVCAN
uFNGlRZPc7Q5JfyNw+OAMb3gLmF2gNyYzguQkWM4sCVDXulIXnNDzl81myTtyJ+hE2MsgffawJ4h
2PhL6H5tqsoxj+VBNLn77wZEF2J96paMAO4GW5nA0yaUp5DbtHxDnCBgLTMuX8zAtNsK9t6kP5ax
cJP2XpvVDz1UNoXZn4Rrbcct3Tt1xjJOTEZEyCLmo1acWs3WS08FJcJJ8C/V0J1FfJmpKf7O6ex3
vBZhUff6YpI+1qKeTx05pJEVGB/+xKPXWcu4Nj+oqr4bxolArwOenQfJ2+kAa0ABwWnkz8dGOi4b
xPc2DKu7vRvjRmYjUR27FkcnuA5hbBp//RgAkLYvXpFdRGi6G7qKsBEoayAR8N5Lh1QLbh8+a6hk
+9exSohOf19T9FIAtVvKsgNyUpqSqDZcg9bsDxw1WeyfXIpuT3KwglIjEbTs+dDxFuWtaJjphz6o
8EYUSuMSyl1Fnss/iV/IISmDjERijjRfjQ9taTezpfAzSwx1Bv9mh8DL/wF+joBPRV/hjSNtX932
nwoalAGS1u5qwF2IGUkCACJUrHcaPNXLvMlPVaJKrJPu4KV1Zij/4Qhvuq/LEvKn7hJlHjz0neQV
ei493ppyXsJoYac2jBgEHOtTE8SUXQH2QnKQSxu0UpcY1CfNrLb81jsRjWGHogN/1mxWzH9hUHta
uChqqf5yg8EtY0JaNjz+O8+fmEvE9tZhqy6SJMQv6VHIxi0HWBe1QNoYF/8SOgDnCa9CW7JWKXTk
otDZy3+zEC2ZAdnwfudZ8PAJG/bs04ocj/1Bmtv+J+fpW5KH5M2p+FR7qgqHX5J0HgRESt9V2cfg
T70JhPAyCopHw8zsn4HAERlnrLZj/aJiW3Ooe/aSAhKinJNN0DowMewQIWHSmqvoGXswirIUMG9V
Dhi5Dezm3O0fpyT+25YNb69ZdmPDCL7FflfGUdqRb1J6LAKYmsb5YGLZfyBFpUVMpECz63ZsZgRk
4eAnU4R5qZjgQ3SJdnzyN5GaxtZ94M7Gv6jVsKWWKJVIISZ+dzPPfN1gcfDpxD43h2flsJDHo+KD
uugEr4EjBBJOecIdrSBo19uh/Z0MA26SpF3tklhIwzUN5EGn7SyT21XMfyXrEv5o7tP52LZwrqJI
z6pQJBPTfnSx8YgsUbGSgG6hH2yCXEwkOTtr3gMU1eEoFyVPiMkhgEF2N8Rivxfj6qb/403jLyQ/
W2CEj1PtssZrk+pox7Lyi9XHGD3icWicuLcd64yvp1hyCPGjVGWkME9GFVRXFWd+exYgOrEQHnXs
L7nOmw61jPgtTPR0NEDgsuGLhUvQiZRZhRKAmuI9l2LgcdYCFPAZL+jkZdIZ8clnF/ZDGdBoZcjj
3AXkyWOh4FHF864EkdUYzAvDLysZ2o4cNO8efJzBraRp/rPJ55RgdjajGSOlsAY/bS6MP0HrvQuy
PEo+H9NnKtH/QxrMUAMpS8+3sQQAIm+VwdW9z+jFt9/rejIlBcK8QPiLkN9wQygU2fs4+YlQpjTo
u5BtCb18bxwCwmuTg0OUPxRz0msc1oDkKD6eyqvZcWhfw1R8BlkxEFZxC6rGq6VUXmwhC6zfy+mh
laDePI00orLMCWAsLpgjXCAnk5enQ8h8HDnIi94uqgPqbiVi9AiLHzgVj0JlZVGn/FL47cmXI66p
v7TPxH9ZPeRIai7EVkycWmVh3H/XKdc5q1cqlA8s0Elj3yGxjYK9C9PrXehQHc/L7Ug+QHKc7l5M
Zw2bWp3sCiZo//a0JjuFR/CQUorg2WSzZEgCoA3SYfiIRPqr0nm2x0aGs+uVrxuduNQfDJ3PloQ1
pw+rcV5TgcfWol4BkL709bNYGhr1tZBQWZsTK+/oYTwqMYOUHncm4we8N+W0Hl+eBpg6IuYapGTf
m88N4TOIc3A4lsc6Uuy28qTEzegRuyOOq0by7akfD5mc0DOMzDm4NivRHs5LkretaWcVEBAoWzTn
Cjl7RQTNeBCjSkoHcztX9jOUGG66zY5BZi3RfAvKQftnzK6fGXdA+gBGk+5pCNn6ekx1Ycjv2rbD
Dn/qo2YdMiyXdblUcuyfyMoO1gUmOxm/J3WEWAUgzu7yDy7tc22hc/Smvd0H/fVEq32KOlbU1uh5
ki57PbWkhD0vW6ZUgMJmn3rCqEl7KU27Eh+CUssCxAxDbmb5F2g10wq0eG7VvryVtRrUHhGjMk65
ybejNEOrrKjCRDl5t93QfY+XA2rCUlRvhfL0MEFYn45QmYleOoq4esbGKbbPqIkmPK/TQEJTlNK6
18WCA4fBCiOwk72dlf1UMQbjFGnWREwnUhMcaOzOo3T/hW90crskI8sWPZUVRrFrF8NBCPFZwYau
qIljiXJXRsh4LJi9eBsoiLO3pTOtdaOSmkyml/h4ik5Qq7f4M9wQN+8QGFh+q3D0WvcpYME6D2+I
EtWAIBzoA8vx/44pTbvYhHakF5xPRp9k1AOvnbf2D2OPf/TNAc2utNwUkmXjuaCr5jZanaO+bLwN
SIHkZv5p9GEu3lHpDPxGsO7mKCDSHWmJh1AXhOxpGbFnMPKQe3YDwI9slNkwUDIxQs3wj5YB1hGy
gmE0kMF75gmejVDZiH4J5IivsDyMRFH7SY6wdxGo29KJ6XV3sZ6Lw5GS5VzvswIKF3tuj4lJhMEG
vTS2LG1uoQLGWs+K++vvGMyuIK8BhVI6TExy67nYiLdK5NMKVFkfmt3OdcI6GI+fBMPUlJb5/Xjk
amSKBR7OgHAMpImlIunmLaEgKQqowwvNsHBhq8mS/qLQm3J0+pdk9wdIl8ToNW2vaXnA4khyUxWs
s3PcPITTJvF0gGYvoBXbaEhGfV66aNhdM9o6lM0M05LxRQUMlqX94kOJwgrpEi59SB8BGJV9sgqK
DtwAoZPNs/vxQtmaBHgVBxlUr1NKMG1ZrBJ8AgAYPeCgK0TGGCYwgEs7CUIhDnBYqaZ1Oiuj7ZB/
M9OA4wchSQ9dBVyI0/drxJjDg2OXfTm/n9AzO8skRGRj8coGpugntBh+KH7BubnRPG35/zO5d9wt
1HIp8zZjMxMCTTtRuCrcmHL97pECbFua02eWBJ7eOrRntTPAZ3xKjnZ0iPUY8bxjkP1y79skKAMh
w49fEiqU2Mj/EDDUBq10i0b/oL2GPFoNdCGbjbaFko8vrT9INJIP9xODANkuIpF4Vu3djtXuVHOJ
tQfXvWunVSUOPuv0VfSwtghJbEI5KmsLrmA10yv4lMAn+88eT4JglMgItaUmC64gnaAHmDDl7Vo8
T392K6txvoChSLkmXKttT20TIXDTftDdLiVtzZeTafZEQ4lmFvEgcuOs3IZpPkfaiMFTHVAKxPMe
VXhwCbVex8LmbVbP9tASdYv7/XLysBYX2VOCB0d9XNDwWFBTIP0sE6bg76ddaawWKuvYH/sEgbV5
/VwXJLIfYy2nRx+Wn2/ok/SjenaagtWyiGUbzBL/FbEMJw/AJO7BngB9zYu4ysWOI9yznOVzEaxn
KRBEjTzpyhmG666X0ppCtzFsYhdlzcvDfwDMOKFl3L3XPEhsBSZAaQ09h2WhEfgcPF12Cai1PMjJ
lI/In0WRLfkM+SKtClN5OcZqx9QhQgE010Hb+RrhIyv4aLWBygQfXQcGgXzjuqPeIwR2H4u74OYB
8gqfway0lcONuH/wSXlLFTrWNgLNtADj8YWALdcmsAMh6PK7Tm2bWKEyO83CpsEfwwCl8IWji74x
OcZn5zIMxA6pGCQjnflekA+t8WNyCfWGVdpAleku4zCLtYW51I254ZkfzEqeEDloq3VTQ8kKM8Ap
cavbuClSgKSG5MlIBCO9P+i8WBUETkvAUT/byXxOc/HSb8LqAUEng2dxQUVmDD5w6tEsgYzpDIV4
i2alYHLMTQBjTrm/Eaa22DdoFxfZLIwNkFnEn6j9eSzOOy5cKpA5DKodTw1zQReo9w6DrdenJN5N
bEQb3i+Wx/LcnpQDlM8IiZgsKaFcc0aVe6pnmuRfM4Qi4WHU5y1AucpnnDqVZzy96TxOz8S/7dqU
mFxcMYdxpi5jtQnYeXi/bFeGwnLLHB4zW29v+GqG8fJaEJvQ86X9RDcz6oa346YOtA3wJAWQUX7c
esNIw1/MckxsSI4QUkQkoF2bUCrcRusaM32XZWeKiW31wY6k40xoNnddBCpfRMULsEbExBvPHfdG
r76tV3uA3EZlRfweXgknz7qIUKNI8iLi7U3b1LI9m4VXTyDKWpaPCcjIIiospiz9EevSEGs8QJ6I
AWqYfmjJVfurw4bgg4L7ok0xJ1WjwM9iNMpy54816kgNF8vwSJxzPGfeXyjm+s5bZ2dCX/Q9TZ/9
5jgLCrPrnbNR8bnCfYOH1wRY4ce8b+WP2far5VMbmjmTfzvanu7YVAW9nByo433EZkGlUIn6u7S5
T47xVT3NZDJ2i5gVY3J+83bt9rZJbE/BgN18ACJaTayOAkKziHSFnUFUehyEnE4yKX3ugXDIxgIg
cAnDr/oNNJTnjLAvYosSNbTwSJNLhT/OD58iSrI+gvq1achwUp6zpewPBNUqKDsCoD0cc3Z3OqD3
n8Gw+6xAubCuEepsvdUyrdL/9KLfBb7jCj3BdbD7Q1cwlLA9mpO2gywgezxR73rcYeNRSwJPvtVB
nXlJJSXHQmWmOzTGoVuc319+IhTwvPhFH55JL62a+FjcV8nAnRsqg+s5/D5qw8cmpCCaWgwFTWx5
wl6QmW4K79WDX2LyqldRcvPgVISZ+awxM9Bl76r5ar9NSDzdODjrAJuXpUzD4oGayK8CuQ1BES4y
6q1S7ZnTaB71K1HHhF93r014sBCNp2liio4Q7UDkr0XeCZJdf13ar+eFfJ21r2lGZEE0kTPgIozZ
7csVWk9529F7LCpoCj5zGUA2NR0WEI0uDqnCOUDCntNZuuUMpQbsOw42fuv3qIBh1SSQosaK2lcC
6oPMdAe9+jnzMHNaUCnJF/UZJrs6ucPsGb0+qpdRMX/1tZTa5RJ6aCHnAbkfo+xK8iobXzUHOPlc
QVsjMK+88KgxW4ACkdmWsdAkCroGgcuQaHcikJQLkeE5bf+w+iIPJ4VRqC2B6s8rjgLAlFkNnoen
Yqvc0QV2dFajt6IWVLPjB3vBd1pQc4TGdGD6h6OWKbFyOLO3qajBhxKclNQTObpW7yKdw3YxBqPQ
EOZJWw2WuAjqNzgFvoVLOQvoXYm9QEBCT+Jz7/ZJIk+9pXlgj0YQLPhsKD6GtKjVEsJM757SRS/v
zTNL0/R1B7x1Qqm2e+MjO1qBT2DLrzI2NkYR5289DRXq+O163UjSvd1XFug9hC+cAP3tmI2H6sEp
LF+gd0sajTWs9NyZmaP3DEuIcXQumzkqa+QlG/jeEUMu2kKRc3KzvnhUw1MuXySO7cyp5yvLTsEn
/JpenNzkY99r+yh/Ql9prhYl1/xI6o9oWjy9WJNdfmp3ojIZMv41DXTvIEB+soOsr+3wO9tkSInP
YYshJwlQLfnA2cxr84hyy51WV5p+psrEJrwv2E01CmvKYzJaLrSX4CRrfp6kc/Nmfhq5a3/KR4Yt
a0y/JE3k7pYt5kLJaDFCVbhbc1MQys4cCoyDm0l5V3gMJyqZOVlAnVy1fIGLBzl+Asqkz1jicR50
lz1jgb7zmNFpk/Fvai9yk8MrJsBhnkz2GNkYCQ01yVkObsMo9cx6yTmgS6TApx6YZ0omFRJ25KWL
vzcozRFciaH8vCD3X3O5fT4SWfqvRTlFscUzAhe7+eKG740FL3HIUvzgDbyOaFz+K29tXO8uIf5D
cI9Hsz2D1ZvRt/HnZnqWZLbzaY6BMqKfBlZSh8Kdcm8AynjE1v8CzRs/GidNOiHqk6rO5ykzRoF9
urELtHvpor8z8DHdPUmmN5l7hdWD+fH43/FcKYdrX3RPCdyiHqMT+KekFBsoa/52Yn8oRu/373Jh
9QXPNAT2KblCc6ThR+1wBZxDAvWlucDlwQG9HJWLjddlK2452kKkfOnnOIV5bgN4fuHDgi4Ou90s
xxHFFp9YPrTszhENotC7edp/1QS0WFHaKWM4v5uDmLtM3ODS3po67nGeQtpNul0r4FGk93lsxs10
OKEzaGLBTUBb+bZhY+LCoG5mE4qeT54YsY1hN7WSjc5V7KVBVQX/7hCVxOFcg4y4sqo8u+YIJX/H
t1fRvsDNdwy3z9RvbrSThmmdGftPM89Zg7qR/Lf3MpnZ9Pym7ujEzlRBjX1ie9OYGD2Wam5rIXEU
cIbAHG1QPQl8YV0BMLtHDW/z2CAMYXRzgQbIl3RcIRg7Do4o/cflRgRX698CYkK8LZzTDR5pqJUd
9CmOC11bxrpo6U0JZl61cKqhNOkHUCMnZ7Y0Vlf8IJXYAGiP14DRFhkJAkZyUdkia5juoqWO4WmL
RNUzkgD8K5PR2AIYt7LfKG6f6O47Tph0vtbUQbqQrMhoSvRPQelsK1oqUFrSPTRYWd6vL3VGNkxY
5CqsvSgStIbId+t67UMe58WPNafZ1wg2AixfiSk3pI8PHcxj01VMPdf8cOPMX603MQL4FNoK/++K
T9fB65nkPDteFM3QuFDl78FznS7yD1HujN4QPoGVhX7lh0w5g1adsTAdA2RpUrbg63/XV6bx31N1
PCwLbfdwhvYsubqaP2Q1wDi+XPpgcueRdrkVMM1D7uRGleQY12zIJMLASysZRTzj2nYHVQvmB1iZ
MBFn8TsO5I8mnFPkMLiJ0pw2wH4JrMR8FfGSh/IiKVQQZ+opeFYNhqiRiF5Gmps0ZXHkDjnBIcjD
5Z6a1irRmc35RSm4j/soACgQDKFa9qT4kAvXVk7m8ZoWLUIlGDNWkgOB1MNTWmb2Psh603VV/hKy
ySHyX1wIvnT7bukmFjzueeoKLs7OP8hKBPFWj/XAOVraNxWY0/5AJ+8LSAtOSt+tMdpdMaHyGtcN
sA2LDNM53QBoDEge285GXO1L8/wDg6T7sCYV61WVbb1rnjimoGCwwjwSA19nvJ05crQYcgAS7UTC
AWk6JX/lcLtrVdm8lAT14lrofNyexxCRMhkOXJXoDTXm0wRgS2NBsrGxJ3MQdOJwPeJX64fCHBGy
3ua7TLmRUxmnTdbsPwG+Br7x0tvCMzawknIu2W8U2QUrT47x7PaTn5nu9k3eNRe1M7rFBJSnVbiR
npS4SaEPkNUdjwJumeFnjv2ArBdDbpgncKILC9VDdvkfN9wFEP/k9YIs88IQOAN/l1UtpCMmLgGJ
eWYw3cuis+tERoKEnGqdpvKMVKSJqk7H54bm9VggsiwCIN57QV2fLi8nszaHderERsGFRkvxn5mi
yDUHMgGvk0TssOe6K2+3UReCd0myHq4DKjXarUqmIVCNUtw989xMLknBtLukM8LRaYtA4f06p1E0
y4R5GVUp/ylt77gA69HvNdeLuLAhm8LkCeNWcky7SOHVeLiPYqAAIXSjNjtTYNgVYpRa0+w/5tXK
afREqLrPY8KK9nYt1gn060sivY57WD2660Zu+A2wRb2sm1I6/2LheoBjQhBFrVeLx4e2YdYtCNcV
PfBdRCrJyIYXCPhPiTQD0KRBDlNwrN1SqdbQnyCNj7aFSKJx5QtmKFWBSH92B/Bae6xdtbxEOT3X
M9j+lNwUsr0ZwCUXR8rvRDB7QzCf4Wq6f3V+AKtBf62bM8k9tmOwTTw7wHs5gArlw6T6VSxCjQAp
G1JdIMVBTA4bA0IWtOvutyWnarymsd0xyIrIBK1C2SNXD73nl2wLxXf0q9lOaeNUWyZ7NY3lI9Nf
Snd+DihgEpiEOncMkPT/ZYkQ73ONVqEaGm9OrGR1Vk5T8/+khZoCa/z+FitG50uzjXDP4bUkuOJC
BUZNq1JK1+DhTfCcyKWw/S4U2pRxiisLxz+SWLfMrb4PZqm1fwjjqT9UACksmGpWt6qJZXbkaC5S
jUQUX8n0buTJEFSi0iFvZiDbiAlxDL3T3EuOcGYYqSgumSoT2GZhgsVAsoKc/BM8S/bcwe6gwSgk
FEvGzG8SDIe5KiOH9UJXxmuXyIxZST9R2cAxWrZM10pG7L+WHARzcR26rO00aVCZQb+r6MVjKSuV
DZBSeul0bZKML8NM4Kdp153mJwtnC6YIbJWkbaLoo1y5U1KaYqX5RGhyfkMe7xfSq6smdEgC3xxG
agdzurOy2IVAC7qSnbPerHOUCXhpZ925E3rAxNqA8Alwur31hFpuv+fmGCI37SawM+GsCRG1iHKy
UJ+N3DOUyqjZtA6bmus2WS/x3UGQhzxy42hgwohMQ4SmYkkE8OOfU6u0ItVUhAII9tM0aUSPV+xI
e3OWvhY2xrChlmvovLFCW8UEDFnj4TOHlI+OJOSduoa86PMA0hYBEw5GWTHHH3R+bnrlqdWhEnCB
SGBtXfK/mGxtHecpoLfZIwISYTEmEDZOJUJgKde2fw/uEqia3fN0DJ3hplJB1cBBVO4enuOo22Yc
JPqlnUUQt0AGrg6lYDdhP4TZU+js8br8sDcOZ/lov9CoXCsEtZuruz+fsad+bPXhicTjB5ym0QdP
agxiqquKD2TaDz71AZfHpgYhVvMy74xwaPRK2JRkD9TER8BepY3U3RwLfvChxFNVyLnGNWabnObV
u5fI/Er/p3S0DsLUr4YSBeMOtfXxExzcurkNsI70C0gMxCv145jSKCjk5BCZOWte8gg3Rpy6VVjF
6Uw/PymLz/i1NokyAaILsrFyrXiO+PjWx1c+km3v86d6NpBJlsr3vei6DzCxGKAp0ogtEYd2zwu2
3e9C/+7Axii9jHDVXJHYojZ4g2mJHkcXx6ZxSZXTiT/C0lL99+9XBIo1w2llP3oWfRQwMTmA+gnv
Pzp6PN5NX+D+pLbXCqIq50bPIPpqfv/Dw395vCr+U6dct3JP3GsME3XFgohuwpTTDupWVDXLt1zq
vrJqTAgZLUOQS7QLOwuZA0MarOZAfwrD0Kdbprh6P+oJzggxvP+OdZvEfmZtSvlH8XQEPm94N1Z/
EjnoU+rpgDqoOr4islwzQaj5WRNZ/ENHNJN7Gk+azJxfcmwdNzdXtMTvPvRm6t5vn78o5OkichKW
NUlan/Fe5m1wnL2KLp/dk0Q/XVRO0Q8K8+aaO03Pl7Wy6gABQBXUabL4f5SCNUMHGq3elkfdM5vB
ZenppHSrLo7rnLbzSQWwNAKF7dbPzEI8kbWhtxj36P1wCpTmfHa0pC65MA5KqCqhbz0OeEf0RPh7
FD7uX6AHYlCXpi3HnhHAUWo7TOcTHz3rVqvGci+xu5b/VQNIzohrT1B+mS94oOIOPmJOXF0Q/938
s15njIyA1ZXddQYhPsmMZV1N/0nqap3Mzfo52yquPccK3g8GNnQ+RsD5ANsgv66/3Qn/UWeRNItc
drjyAz8Q50V5SVkl3hSpIaAz3aClIeR2QmvvKJARyRgt4nveQ8Bjrmi13Azj5AI8KXdgjxv3a8sQ
gn+OQwFLzhE7omVXybsssqoHpXYrtAaJEoz4P2KSe/KVHQquzHwFUwxI+ig38rSPTnqbOkxxEV0U
X92PoeTj78LzVQ3RCGE7Tj7B8qPRw4uCLMxMzO6ZIVK4vPBqK0xXgMmE9q9cleq9+ntqK2GxLsaN
ERzhZKTUPSFriaNjX66jxqk7q7VZJPoDGIQe5Z3I7ZGqFT5OrBmtpCRYDlnwptKD6n85CiQEr2DB
DIFG7SA5iv0IQSGqxYGgzBhNAhmp+2Gy9TsbsglD1FbfEzpWkZi1l8T/0UaciOeiA0GTtaanF2vH
RldNoV2YJcd7W6xrPC0a4ETndGz9r+nFCuzGtJsmPCmakkvCGLV6tP9HtjaUcd0LnnbTXOdKn6RR
qwgcNRAcwWz8PktpuXXrTVOnsG0LZUgaEHaUNE5YNNV0/Q+QjIfLEDsYGdB8O0pSCx/FqQM1Z0H/
bwI9Hy+wQMQKdV2m4KxLWR8eLrvji7NUEprGmSiN18zvNl5R6Gk6RaE4i+bR4bkJ2f/GAktz3CGk
PQ9XzyRre8sxCo7TIEj5zlqBwunA73+0xF/O6MgD63VpefIV7aClTcWChF1kxf6t5NXLDZmRQTL2
O/gUbi3lj3hvcfyU/tX5hVrfFKFi2O7GAgCI+rZBQmXKRDYEqtnoORd60Foaf+JxYiW7AP4+K2+o
/xgBIU92EsaiN2lH84qEcRfTW4+s3Jo80flZXuO7KwngmrsEah7xJcDTxcRa1TQ7AEt1Z5+6P407
rwO0UDom3AkIGtZ+0QQ1iBL9mJ+aJa+MBvV+UmkRNDWuqJLq2QhhktYVzmZ+yiOfmk9hzT1X1/Rq
AS64lv713uTRaOuOSoH2E064TPNav/K78WISBD970lz/hC0qSVU7wEqS60SD4WdmqlT02jUHJJq8
8s1aM7b/nFbqRC1KDAvA+yWuVa1YMghZChmGFOlFdJPoWPpHRhqBS6bGK6blno10MgSOmwzZbBYk
OLbHGvTG7lfOdazjotZubf+Qd/+3zbEyvYXQPyv/JSKD/fX/hvvHKhmvS937/1eQ5D6Bk/23oDBu
DRkz+E7km6sre/3Bt3Q9s6lE+nKzyKADIUIuIvKq3weBQ272b9fo53hM8JRcPXulsuaIp0z+yA7A
QUHF7fm9FuB9JwA18/bjtkClnELvTcwjcwS7E/Zx9wfRISvcHHgrIq1IFYHpQWN2uKEXjN5Nn6zf
v30i+Grk4JmC4rhd0v9dUhtESrEddV/aJngYUlBDl35eunKaIvbt5ELfia+xHUe3ec1JSdyhrxZJ
+tvDMOCudrHzldk2ARUFW2VmUbr0rOkpr0vNz/K+mwsXRoJD7vOZyOcCiNhpiN2JsAyKokL+h5QK
e8fiSnv3acHBPW3lEp9j28KK7jvRjmxH0HONBTHUUCeCuk00rXV4faOdkmRykGPdxA0hDgpnDe5X
8hUWd5RPN4iEXeRSb34Dpe3p0oD/3y5DUPhmU453rRqyXlsUGsRXbIMkhuAeEGeO+irxcCDUfqfT
gYK5iE3gtrZibdB1XOddjV2sW6xH30gG+pwXgkpQ7w2/CQSLsHlp4FZ5TK8CXAe0b2gTw1+/XVL+
jRRKwi55Jdw1tKZxBzHwur5ilkUMEnpmVE1Db3TSE7wsTZqn3rcsBOt1iPjgpRTbVfLUHHLaCZxe
XgP9CpSIdEd7MDMhJoo1MMBslHuyi3BmnkQp5pUSPuhvCWgCOl8Gx5HAR3Ren7tY15zy/XYIokXy
zgRNdYAkQNlYoD+1PUxVkMfCYXPOHs8XPCZ+EFUcQr4GLO7ZSAI/em3n2rtaF/8igeNXzv30oonp
z3ci/3tKF13nA1HOr0bQ29HBxffw4eQMgwGINy+qVrqugeIDCzp9fu91vQvQvHpj1z6J2KQ8neQB
MEKayA2VLhh97T8xztoTBf8juEVC+sAvsMyP4bpKVTI4eDgLf2EXhUlT6+/2qQbUH/C1qEDCedaH
iVuoxuDAIMoOC70RguxdnbOiqdQyJ2//Ea4JRemFAqhUfar3MFkNs2Dp7E0qDvvyCIquMCzFsPXM
XLvcviBiOfGuoEcJ94GFgkiKSO9t9snqWHR5YrcgNhno6EGETlP6IDAUmYfDgfmR6ljwMsywKRDs
1e/803fd+OD0OSo6WkMtJTT8seyaj72btHcrp3E9edXuT72+GcuTSNbD2OhP//6NGcbYHO1kn0rS
QsMotwcNXjtvLjtr7fD8qSRa7E5EBuMfVVytG3XJpGgoDjSkJUP//REHuoxkBS4HvPkw9NA38APm
W0SeTcicf7vNxGEZ5xPICptrNY8s/JDJwuADyJlVdr2YaKrtlPqDer14qb2U8x8HL/sxTFcuS6wF
Mcoep/CcesVzTriqUFlCGLmY5jZ0xQOnuPFvN4EWW2rkOz2PBmiIYd5dtoM009amUvbg0lcr6FPh
KBeVjt8s2HW45JCuhDCK8aNkqJsrB+XFNquK35JI80Fa/pHc+yXtRSXm5U/Te4sd7oTj0capbt4Q
042X2srJkAObzGcNH05TsZJJ9F9fDgEMBRaFdbcE+u+9HGXssRSSro3IXf+V+AZgRKhWDxsAhtGJ
Jmh7xWmDlFwZEjgq0AhfxkGm8sM8xIKz4LFsQ2nHRMblUUk5MleNVNV3pN/i5jjE1EPYDN1iovK/
W+FvNIXw3TICZ+HKObtLhBxGyYL8+w2zX8W6XMPMzn25T0roPepo868eO8d5hJ+mJfkmcESc+wPq
Fsx+6hhsfIfoFuxygPKh5FWOvcKbdHT58FYCuUnh+vcIN+eYKZ33f6awcucPki+cOrQfJJkr4u9k
YCRNK7n9fNL7dk31gJxwEY4/YWhjCQkfu56pHb0dTFMD+QoHELZxyhJn/Zu8YoJLT7tVhs6tjkvY
ZbaLQfuZKpVCmiQzOPbkDN1t9Ngh7tIi5/i/HLYIohUMpdybw6odL0t1exjY4G7kr7NlMBppQs+Y
BmXw7pboP0zM8kZVYq50W8mjnDwnDD66iKEL0pxBQWqw6fKx9EO4fEStr+4On/bOecMx3PSV7o9Y
quf6+bahS2C33X9ta6qm+hXVS4RqBO2iFhJyM4puja7M7hdleC0612nShucT06OenCEltB8fR2Nd
CZBP6pdot3CCMBBhaI26FzAS17OWyAcDF1UV/b0bdjWcCZZaN+J/tBUJ2Yx7gaQs6SxpX58t/q9i
tO6Kf1JYgAkkFtBdvA9wUCHzNtJ1k/kRs89LdIiHUHhZuo8AWxDETKKTbNH3Sl+2ptUdfvwKgsRQ
Tfs7IOOoLnym4eXszjXb+SP2FEIDRexE6lBfb0gzum8vfRaIB4dWIKdP3hb6UaRRN3dKBapkuYDv
k1YuVtSvKik62y0fvzd7/cuEiZ1kUujeqHw7etyx8VWaR4Sp3VRudPRcMJDZlCfSLb48NpN1WVDw
1kJLj3pyU0zaRE7oRfWuAh71QFDfftdDAA41Rw5Kg2p+zfm/dI/zdngcP7HHMLRZ1P6te3TXrLdN
avJn8nCapZ98BmZsg5pDZxSzSIsBtI3rOLnWFx7tP9NOaaJXUfIX47ONp3hNLLI/b7FvkOakmod/
pU7+eViOasnamH7D9G6Oiy6XDEd9R3fJxqjPfvltR4Gq8xsVyrqX6lSzYo95HGhpsdMvXI3ULLXL
iZG+sgqlkYIwsOLW1bby+lQ2GSoTPK9kKKXCkn6Q91nyZieNup/KVqWS9ZsDS1Jw7V5HS7nMkQPh
FsrJgI8dWSENkcocljXoCZ2JNlZI7hClSuXsNpi+92cj6mm3Tgt9rv9d5M2ZADSYQ1/oSEzzArLC
ONx140RMJ1R1YqsP01+HnlVtkw61iA8kr/XqNmLgU9WuiFvlvnsWQeF6cVUbZjYpdiuKJKMCru85
30TEzGkZAWVFSeASWUn4eMRsQ32plyN2oY2IAOgRvU4c2cjeJy85GuZ5BdaUWPlHklaRk0/blPRK
8LMoZlFNvpQgoB1RI1Tj7gPfgfYPE3CkqhgR5aKbl0R/sLCuRKm0/p97BWjKGOHabeOkahukckQi
tnxjwyXHrqDrsfd1vCYDScu8QqeNY6Z0SBYJAnPBjEQsKWntQpRheDZS7GfoGMBoEPuYcXTz4jKw
YDXdSLakQvlTzIL/dq4CDBWFDgiHlDq6+k0BG8D+uWnekMxtfXOhSPBzZZEA7vPm92hdQ0LmMvPp
m95eko+1wm4cy2fvrZTr/mmnN88uCgZSXr7SxHzkE7GG+n9OSN16kuzMK2HGnJx7AtkFio7odtIT
5LmGWWjzItWXFdQz+qwwdIVSj78tD5mgXslZat33OsSNhlzva8dK8ad2eK1nNuL+dAA/gdIsIpaj
9AfPaVsai/XxdJBNbVhGyZcZO/Nz3Q5zE9RwXhMSkYEqMz6ugq1MEZzE2Nu0MnF8M5Z/Ttdv8DJP
JjDnKre/lCHzM4dUgjIP2zNTsJLP6oaeCXFF+pzonk6MZx54fFrYFJqkiqFUF0HqJOE3cgNr7bq/
w9RcZqtHqaTPwqJpG/Rc1ZZWQr9r4Sxp6qhd6HEkmG8z+dDfiVxsztDUaKc0KW1SWlDbR16ixtc3
+u7OQyT/EJW9AjvVCV4zwbNfrxA914oYis6amc0Vg8xUc91fd0KOvBAhIGueINnczZmVAA2VtdZh
aq4JKNXyH7uAapMJ0uD0bc3RDxxw9L6WpS78YYrmvaMirajPSc8kNuOGIAAwJJVENhrtwvn3H2hS
EiSb3F7Kh9AQjbc+h62hK3T1tI7VoqZLp09r/6D+MCIZwMOAoV/QLNLewlDtl0tjtDjEvchp++tg
zv+6EHK9bDV70HqKG8h+N40lBQfKu+x+mcuNOXDYCGYlvnyD4G3tLITdwC+xqqb4ATpzPiJRDaDg
Cgid+a+ZzEjLP+/wmoDuiqqoKeoBIXV2yFWkO2ncuMOJoKBHkUvjhsWRyV4ujvTiMMS4Sx1morjB
0Ltjc1xxW/WYKfVkJl1tezPFawNL27IbwepWAZmTFWYsGb88mtY7A7lf6OBLKCoggw6PXDsNRLLX
DHPwBiW93rJ+dYcu5ZBIb/+jRuBMgJmFM/EyH1uQYSfnjMPiIcjGundxnaq1ERUopgzc3OPXbPR5
6vn0n3aCSszWi3ZZRSAjXRcZM+cRRh2xFgAevTUcQ8BdcAFCYLE8/D05CoxG8tMQ7hIGpyo7MvQ9
5zovzJnY3Xm4haRtKgfOj3nnPxrie5TKfZzq+lq5nKaTTMIYZuaRkQaqOmtI882ufdTrAR22htiy
hbP1sg4fe0mQtvOt8KuMzA+z9x2KxW0R7W1nDPP/n+q9fJQY1PDu50q3Fv3J2+6fbFdmqxUAcyxV
nkXtIYwz8Yf0sQd3zw6+nrm7LCGsj1Y1T0jKd4U/jw39pnmVPZrreaUTr5HStgpueBFiT9DjRcjf
CxLwZH7l8JKEGK9CeiH4/Os0ZRf1lz3zR/UjLuONXrUFCUZUuzBBNjIj1+HOuV8QYZjMMs1GVDKK
Zu18wzvFz9kwvqBWFVRZQIu3slV00PFvS98QYBDgIXGtW26tKRIC99CyTBT7rvy6/Nqdl0oyWR8D
WonOuLJzEasSkCqJr9meerAESSi2Mh3E9tNYssxyCTiuVUzCAV2aJYDXny6Dd+l/R2H78nijSIeE
Z+wa7Z3ChUmBGUOI/xKIiw5NTLOMkBo0GHLApMk/K/CHT9r9ftNlyG4FisAcACjhdEPocIZVjuG+
aBrT7c6xV+EcdCBgHsZpyp6Eh6yEuAAF+WSZtm9vVLcirpAnocc0Y7VTAXEFXRhwfhQlKjVu0oQ2
/9nqsVUs4iM8B3oUWqpOvYN5DNX9ufmk8ZJDsc5OUT2LffNkR3ftHGC29hz3h4zXDdC3t1ZA+unU
QssUYyKJuJ+N4f8AvcCiB8tqXfYwG4ZBOuvRVeTCtM4XnrF5KWTJ+8E9IQXlSIK6/BDZBSMN2KUI
KK6AOVdGXQVTm0hfdkw7kmMKFWhsI93jNR8ayRrx5IzbvXm9wCBkDlDLlHwcrYdUUS65z3oBoVHR
Qq3UNty/x5nq7Jt8r3vcp4funVwlfhxsXsmEcx3JWEA6t3pycLdu7HV+ofLtY9eIRs23/84MfZSN
HYd+MRzHDftuwj+2tFPF3pFmLTKFt+HYcg5sAbktk2Fm/CRwVJbkQqGHP/MkeeBpnVxkUs5ad7Xr
f2T0EvJvFkbftyVMFHpthkonnOxqn/9QJIpEvNxmP++Cpl7FB8415letM0GrhtA1R308mz65S93b
/GYf/ArTfUf+saq7RpwXtR3ks68hmK9ljVsbLBcnr/SkLxwgL+WWsSsEwpWNPNp/KCp8p49LCEkB
zMYJj13rsnAqUFDabrgpmQrN/s1LXu4kj7t0tZCOZ9pec1r8qaThkbZJ3xTyrtIkaprZ4BT3GxTO
z7cKMuaDubZdKge5wiORfUDehEyP3626A6HVNBPGVchDWMZjrlcWVPqDfLrVWTcYe0GaqgQgRF6f
qvqzAOPkqtDnyvhhRIO2OA90B1Bw5Rm7FymjbBuxWwj4bcMxzfmSvnIN/oec2E6FJaOGtvwLO6JG
YMa+ByEpe5u+ZBwljjcIma08c2DKA9Vor7y/uL/oQGYQaCtKdDojjKOgmiPPrOfV3FvJNkDp308F
4ZsuDd1ZRYL2rZadOSEDAfKWNW8d3Fct8tUMUSdhSNpayXTCZl3F8m5K+L0dhXC0YNGwNrIYZiko
LdEqiZE7xiaK534s+47w8bHBAXGa0FvqPld77z2TRIUtbzpeBHGwcg9DCgAxM8OHRduJ9x9xXVaZ
jAxPWgFN5gM/u2YDgX1Uj4KfYO38eHGuvKeuqJeCk33Zlwg9CKkJtlWnEwrGjJ5h06wkXFqL3vYM
YQqbybhFWLHKZVCMIunScVNNjR4TLUKbMCx860dhxR93I+WXBzFOGf79Giv9jlQXwv4mz+jPY16Q
svktiq5U2qFtxGWatDVQmLlVN0Cdval2YwaBlrdDAzSniWAXhD6nzJLjAJPxAmsAOOof9UIsFvWM
aNTEqfzNwof65gLgkwljVHVe+xYL4zYQfz58EAhMRm271E67rPdLnqPJwiXAlb3pr2F5Qgnc5ytF
nXeZQ1yc3FQ2CUB5zbMir5jEVrxS+Lv3gGSRskuL2mwU3cj48ogoCO+seI8K58So3NdbYcIi7/N8
CE3kp6mQ1K4WCMYXad//3jMlyZMmqgL5wT29LU9CIL8pooyqHPyBkE0qKqjdKFEwyD6s8z2qiw3q
wq42eDkr96g1Mb+Cpe7HCh3Ml/qO+8nRgcrJoX7XatvxZQhTZjPbB0jCNU+mdlIsl8/d5uLBS78u
K5+1FCKkvA0Om45EPb42k4NzUE/iGMop3XQ1TYmXduDvfL+MFEDwCq4amYxwhWOAQ51GukErBRpm
Fjml36lKMDeKl6KmEOsrx1RBNeKLCmNKWLBpl4cE2U621wNo6GHQVR3yqgBgPtZ6RofmREGmy8Wg
PcOHOleNaNDixzUzmsXusaMlh0Hog5BIhYutDqw6ZrRXLVywaZBPqPWAnw8vrvK6bYTzK8xgb6Ai
OpGYL+SlgHncln8Zf0EO6ZVhdlXCZBvyG2TrliUvz5UEyLAWlPyRJKxC5z0fUGfL2omEz0f/mdND
LGnaa9fA0NKVAR+cutvu/e+wytLCKZTrAeAgKPLASr3WiE1yk5gik/NQir3IDueYrdOWaf+DOxOQ
GXmcZuLZ5IU/WVgnqkW2PVknoQopb1ctqBUrQmggIhw7+6wCr7IMPfcQpNCSbp47EF5S4J3y3ub8
pP6utIFU0YVC11ZC9dR557PoH+Dma/KB/dFppf60KQje5RIvLZtF+lSWtgNgyeP3O1B/ARV0kj/8
pI8WiTbSKEBLAiky/2BFDgtmk9ayIVD/hYU1+lY50oBWlr39TlnGhXTcvyy1r5TU5vMnNTLpqmmN
b/+H9srCNo8/aaQlcizpnB5/9uiqRsHpXj8gRLNnCY20vnzXXYB2DI0f4X+FQSLb5DR7oA47SZF3
aZg1w6z8WD5BhPiCk9eQTUqJta+5m+qdGlkpiaYywTE2OVKgwCl8ioX0JM2dSHEeTligYxyBK9Zl
pSkNJ+CPLY8zo2c/5rKK/qrsavy+3zKSTCCODj2VMTgzQZ2DibpJa+xgaQp7ouWJs0n+6kWSG7oL
HQPOv0x/XB6ywUcwb3ujHvFI9ubBlYAWK2RGGgm9PGQzHF8hXcUXHI9L+5ef1AMSQZt7cZsOmGkW
dAtJhvSXXUXx+jWfOtTsceCEdG/Ewew5pwrPoRrVmewQdHvR3qP0Q5jPOTQ2iDFbOHjQSYlugr63
Mkuxs119bczs/mrwD0bG+n7Q7p59tuyEXVdmtj5ApXwlknB00VjBMoCF1eEw9M9ocheI+bo0JLKW
MC/grGBXwJc2LXV13Onocz14HpJStFBGP1KA9B1yP3N9x4co9EalTTbGtOcsMnuHZrWoANmhkJob
mFO7WKLnDmBDDZDyd9WkjBavN+Ik7uc42TBXxffUaJsFnnKQFsVh8kL2txvFfltzyEFNZDvRe5m1
HqAtbKkOd3JrYfVUd2nP/Swb0TlNg8wKHno+YHjjYG3ISNC4nQgLau+JC+FMKlwLZK+p2mv2fAri
fNmu2hXiFcTfe7OboIzhje1beOkhkGf9EIonzDQwIkMxOl97L1Uo2ZHJWucpha1+hDWfXNqIDrGu
gA+mORUeacXGNJDnYSXrwECUTXkiY55kaYVD4G+kjPp9v1LudvvHdGeR60jqQYrkFbf1L6mic2th
ooqJI19YUTMv/yNfUW0FaBaazprWushWz+xZOvCFwTKnkkt13RhsKSEn2j2LDfWeemsmq7wxtUci
bg1/LtBbZLBK6pRTfxe5dcc4lwMY8hm9yaWMECMqoKOjPam+xW83+NiRqiU1PLzglCReIdWrpkZ0
QuGAKQB1IKWWqiG2j6D6fLHiCcupndnf0LjG96YQGpzUrCghYmBcC2RjRANTdRwkH6yBIOkgthQA
rybhOQYfOTKUr+LsA7HmvFjcNh0WqglyioWqCMWuPddzc9jlLRUEKpPxTZXuujxKafs1IFJvsipM
O/WcRZocaSzKpxDBuJc/ozttzOJJ6yFSGfRKzKSc7tR1NW89tdVJYjDrRz/2BIADoC12diz4A55z
0JSJJ81c0jwzEaN0BMmJbhXA0pcaV929lsdIHX73JXubXMGREbvd3keX4aZNjOdB0e+3Fxb0WgNt
3sasEpz6ShACNHq/DOV2gO7v9sz3clyI4QJYyUo1SJsd2426kyuLI8aYLoOWtGzL/5hfXCPjtuOc
rVrV627R7KsNtc+98GgXmkUjukQDkucgH0mT6YDko68iCpV/QQdzExDkxgsoyEhsks1jXedo9a9s
ui2PtWY+f14KuLn9rty65Bsn+w12g858wcFI/r4QxhL64Fbl0Ie10rzgS1POMyobu4pxvFZAdE5D
Kth3BA/8XpF/uNqWpv7uUNju8q9tQz9PuMk2+m46LKriKsfWHEWc0TWRRuadQasv9yc4Gcg3ry5a
WqaV/OHkKOmXbfHwJ6bTJud+WdHr9P2VT5R3/v/FgnNrgBJq/wc2SaRVepdadrClE1lt5GcFc2IU
rdca9oKfjl7PRA4o7HOfVGz4Cer7M5D38wYAdfxq907M/qiecXv0cLDvuK42uQopNm0yI/ncTHUN
1HN1RZfZpFaLv39C64ysTe4kPRuABkTIMV7eWqppg1hRJ8wBxcAbeYT4CmlAwlc7RG1HfSX5Wdu5
EvTBrKI2WVUjYxnfZPlqoPcp+rY+1V6rbBA4w1zhQduUrYIzD9mBxlC+7CjIppaV0fqB8uhUSLI0
4WVlvtBQ7yS440Z+TLBzPUHMtPYR+tiEhwgQLBk1ZgdPwT8yoBh5lxeuNIalrI8x67Qyj6rVR+4Y
8DZrEX8t9qXkrFEzjtqEVJmpgOjcSVvPIv2Bfu2gVxts8CvavU6vLJSannPjJlAUZ12IaZL3bmfZ
FYgs5DAJPXpKR36h1euGTolmrm+U9k3ua/qdwUqjLumHwAzTIU1H98a5W25BMltJgmHV5gUV5VD1
Umv0DC1FQZ9tdCqYST7QllsmR8TYFiFA/20JMdO4X4k2KPmGkTQEnWzsh5lVvChVR4zxxe2jACDY
ZiCAFI7wa6R7MqWfuwFNi09GlM1MuG+ujbgIXx4lCSpWkRjWAIu8yzngE/19IQMVVU9e0o8Sedzc
OXJF9h5BfAMcJa37ZVwqB2UK/IzgbQILq/vxStMWRZTygw4mhWzsgG6ZS8ChsZt0YyBKZRKzmbLK
mQu99bqJ1DK2dPJ5Na/BJgu/JJQLAzozEIusIOSC0M6Qsv0/k5N64Jw45/u8Jsnf0ZkGoQYPbg7F
Sv71CC2D1mLNac1wvUPlN7bhnNHrI8JmxGZU01TrUBv83EQIp2nnGiESEwY38Fq7bnO733P92JG0
dFpR1fAjUC1+nVSSes7bXTurqwTLnav5VfADMRPfYC6koBtIaG420wr+LBJeYoPt5shMkZajkJXs
cl9fJh9uqKNKOGJC8Rg79a25/P+FIy05JR71WJaJGf9c/JNsvVtSWn8TbWzv3dEwBr2IRi9crLiL
gfNNLbALyxKIOIlaBo1LUAqQLhArBr2VRLKjAa9JFeHcQTzCCTvnZ8nSKeHFyFY2TZb+BDgeQrwS
zv7y0TuqO2606lOv+nI7NZ9OP7ZaXRN4+WwrbUlOC5BPNe+qImzPm9d2MGSd1OotsN4F4w8Jl1RO
Bpjm2Yu6/cwYxTwRWJ8H4ubIcWFd25U/tc5K/I98GSQ7nGUDxSodKdy95bhStw7KldLkxQSDYut6
VXP0IBuIZ5uAPxtVbzH2niyWaXOF7nUejOFCoQD1b7SOJ7IClG7r4wPQB8XkUARlAOUG8MhtM04f
M7fxwBRhWzMnYOYxI0pIOLhK50t2Uwpp81plBQSh+PYlHxJYa3hjaCx2gLDn9KcttTHuiAROL7Kb
nwf22yilhPWT007c3sfUDVkKEWDR20L4kJmm0IzVD5uEs8QVVeiiYrXSz5ctGGaCRfkNiXIcGpbl
MMJEumhN+4IUYCc6D8RJk8MOYh6kY294FlRuTvsBeGH6V4RkoyDrH1d6Ed2tvi2rdCWPBylEtcmq
QPHDnNplVxkA+z24fh0MvLQHJJik6XesAm2c5SWX1A7BXOCe1USDufI/ojYAFrylC84alpV1aPdm
nILGouomVRcoTqlZUmNhgGpwZxCw8/o93Jvt1+daAwJ0glA+4w5dP7c6X7yJOoCu51w/WnbtMXaO
u0H5e7tUFmFUyc5uk9FF+Ox7Wq9E2bGUCuuP/SprR0EPN9V8ATaAyqhV/GJk2OXPXYMjuqpySqTq
kPvO08ic9qj9CNcuFnQhzcf02m7r4WXykM8nt2QvgFB54TLwuKouiQGjSzYng4+gFTCcRxdZRbns
YdAUqGrdcBO6V2fo+HkR1qbJP4BuDKeYmp9efSdZr9tTDgIatCBdhyB7f+MFA8/PhUW0yBjX/yFu
YTCTw1uh66bPMuF5AKvWTguDbtm2DP0yBfLsrQJk7lTFfKpfWmpGOmKrlH56skYd2YXBFCkLv6o9
3VxhKd1m5Q/FgmvnFVgfsml5KRea8EZ9dgcKDeliu3LhhxW90BN00o858IaUFj/coP7eUQ6IBgmM
MMujJgrm/RP48vRLCx8qjMJCjrSUQgp6z+onwKp62qXmLLyTrEuQzUMxmcb0e7PqDWdIVRzGIHU/
f4Ur/w9z7wAoIkEA5K7Ob17NIVgiNOwQGNps+zmA8d9JElykfF5xMitNyenZfC16m6kqiYPPrYeU
Jytx5/UFe4TNT8yg6W/6NI1pNOryGYCe8M5pOC1PLtgd+VVm31cfqe8741DB/OOurN9bVfyL1gMU
O3qnVyYlNwzJ2YnMoWQPWX/lzLzrJnKRQT78XGLA413FR97jOnMCSgRsNIn0n/dlXcUpvPfGXD/F
LR4basYMIrQZW8u446GW0EeyB8eeaM3A/tJz4aWskRzNziq9KLK2Yk7VWVip0/yPfvmiVbO89a22
2QqtHSGUcAo9HssJIad4y0CwskDv3sT5EJxkXCcCb8Cwcx+Fq5zj6BoZ/lofyhxV5XSrNY2CONkj
KcNcHfR1pkxKwXKcAizIsxXhzvRaJgVgXcp5YyiI+7hc2diyJI63958EzQOi/E23ONzl8NWPB0HZ
mvLoDcmKcBVkanVM9omSJueP8Q09PwnpIdH6FJfAtQGJyYna5JcXDI/KNZvqZH8vn1TR3UL2D/Ci
LMCy16lGpbPij5w40IOaW7aVQAVEf6lLWbfviiTy6y1y2icNQPO0HG3Dcq/8WTnP0RZtZhBeEnQF
vtAbE9N6jChk4D8ZH23ZbYLRjyHent4KajD+MM12lZLeJUP4duxKkhq1+O9NlTZWodF5DrjNU3Ld
JXakoTh1JcghjyJCkcAkOzySJqtYZZm2Y1tOeH8qDJSnxrm/w0pjblDhQ+A7Fbm3cLsyp1fYImqB
1u3ggTC7FJv8PFlLTZGzLH/IAjy/i+j16+IP9ujMM7M1yd2myEb51nvW5Kxf61oG6z+mkfdrk2sf
YM8OdTRmUy3y1t+cMBTiOypSD00SuxqdAL92HmB7mD2yk29Or5iKPyyssasywBMvph1HZZ04t0xm
PHFRdia1sMQ2EEBmwQd22UslHhf0mjS1yyzjKLPVpvIrH+PkMd+bUY3L4fDtHRFXI7KrUulS+d+K
mAnVhj//jlIfRUQJwD03Dd1GpKRriCdxmHwPchdpcPtaizNYwZRh8/6/DW/HH9aChZM2sm2hsaq2
TVLIOkYHCkkrXbgaaUP9u/e7ulEYUl82oQ/5pXIDCUtVgfAs71mO4U2OLLLyiMUUUSF8IA3D+rV6
TwZXOwEjaQeR4iuRrnWPzkVrb8iO9jE9u8JcPQRnEMrBrOux8F4Byg96eDkpwAa4gjgQ1YQNYjoy
N1TC0F6iV/o8wuHWQ2n9fWyd6CERyjXxqGu8l8UdJoT/Ytl2gGXHJr/0lW/uIluubSmrE2c785vo
GnnsSSSQc1a4ZBrdDoT2GgSkDnJ/uM1nZdltchsyBhumwrGH9G1OaKFAOraxV+oac2Qj5nWEc6TL
dy9akpGp0r2DwNvhPRVxhTaknXvGOrQG7Wa5UG8o5BvdrHylj1p/OCugyhmjT222gXF3OSfVm+8k
RK9Zohf2NyNrKjNwIbi2JEpSa5ivl2ba3SiJeEpm8c5Eyv+ksyDN5PPysEjZxTYNU+heCUMr1Kye
pLXkp22LLHUnesgI4oEU/dh36Fyps02LWsGH25XDUnmS3wqoB0F7j/UZ4hIX10CfE1zNjFO5kuVE
sov1anmYcL1lBXskMyk46HcqAA8lbajLAuKQxusHGwzCSzGuZZXe9C58cB9M9b35dOKmP0bRlSrs
4XH+t7QWwV6jZvNh2K3+HNKnntJhLNL42xjslSxLrdDa9CSbvmfuui3ZDzhC7WbM+cwUYl00Knji
tCS4U3ttadwNeWrAk48WNnncaQXNfVIzb/F2OsdlwnlZJSdnD+1BnJTuuqTZLR2dVMdABDKzmYDU
Co9Hyg4l/5vzKXMsLRGbAczrNkiZpzdCPv6f7UYACM1nODt4WrhySKUifV0tZIRjQs1PReSnwb6C
2SPZaAGo1+NYJRjDLIbwk5eiqzwmgqvn2hbgtq04bof2GhTRfAplHO0uzmOJUbWtS09c4pvFsO2x
ViPOGLJHNm3h7DH9jUCQ/lOtgPlcQ1IXjwRAaVokoTJtsddRc0XD/obpZn/WApnEA8hTgZVdpZHO
7wgGVrI2nBytROYagC3Ucjr+Iex7EWyvzc2fs5p2ETMzqOEBU2GoMhNP2CIz0ZEdg64h/yitnBmv
+QHwQ/nBsqAgAWNLuYesL+IfmYVV1c2l0DIBFW1PizqWHGBbliU1xmenLCYBNHmXwpNk2uV49o73
yFtYePEJGQ8OAuGeqD3VP97YCG7pOjfeCuQXxjKfJmEzInGXGzvo3Tks/Q4udSyjhc/IedIYcMo5
vB7M/t6cT3SU5Tmz29mfUrGag0PathYr5IXa5k78o2AfzWMF5l3B968gD+1OjwsgQ2M9k9g+iniq
OwCr+/O/Wv7JZi327U9kLYBEDUOahMDg19zy1t855eUJREVCV7vJ9rdxvhCxYp5aOk6XRw70tf77
NMGn2UG03lObXA+OIHwjXQSazkEZ84wip39o/nbY8e/Butm6VfgJuS2q7j6kgdqhDvgBuaUapmci
AXnJ8CaZi+GFbRI8WnhC897WZjZROCpO+SrAU2aUtBLqhcSAv1yJ89vMN/VePwOBxD5+dKMlBjm9
A4tiGf0r1xMDxfCSZ4ox+U54kVC00n3CFPsUKkBnRJjOVBiXCcYEyYrEg23Sn5QDO5lWHcym0CjG
4IpOltzraT3Y14LCaf3fwR8K4sHB2A3dTru63svwEWKvKi39ZYZ3JSCWXrJw4keoxJg+ZLtm7hhN
kszmzawQ08qTHUm+UU0uwYW5Ri+x0JvBmtjX+To95/pb9+uPg8K47GR7kspymwaaSOmyRM9pkjKi
muIoQsDKqzm9X3YzTwC15HXXY9RdvG8KJylTg3xL8EsZMRoxDTE4Z0YEci0lM5NWW/ZZye4cZ0IF
4l1NL9XCH2mdMFc+XX/0oeycQYHKBB/r8j0wnLiMscMU80tTUqb4M84iRYK3TwNGEepGG0dl3GGM
OjE0T9osl5/UG3aOyu0/+xjLTCbvp6iEBucAR54X6SgifMRkqD9qc6x5M/vJj/7ldnNT2kytWnWv
kJpkIO6ylLM/Ax67VbBAqfmug0GN2REWeSMfe0BtmBNbhVg+rBtLx0EBAZwlojGpfUCPWi6JiIpI
RcBqAG4ziEPMerfN2/t7kmOoq+Ra9UlfLKfY4mlz8mMMP84AmEugoF1QYFGS9MUo+fwN1f2Z7D5c
cMdka5xD+jY/CbK2OHc6WGi1+khI5lbAhiLbyblKvl4odZVG9LU3u9wPWqNzJ2+DmHcj4NoyqxAi
CVh92s18lWBpChJ00ZksvJ6p1LCJlKlggKBQ+v2psm+D3f48mT8wWD3yVJBF6XCE9/CyGopF+Rka
CpXEm/7rJmH/m3dISlVehdef2MlzSu5qD/b6yEPK+LjOSE6m3oqZ7ReCg6OEUQYNNcfmP6gpA+j0
3mGRAM2aO6nm5hRktPkAqy4SO/cZYlF27qJx74g3uBX/lSDoXo0kCU2FKOIqn+UZ6hd9piNpLzan
l6MzHLOGws5o95wSvj5fr3Jxw5ltuMl7dTeBH/KfE+qA2pGzHCWDVidUIgzW3v1rzCGV5Jfeg/Hx
YY16n/25eYPxG3picJgA5JlS5hDo3rvkLl8J9cje5DVWW14lF+G0ZdNc66/SQ9Eid3YzsW5me79p
tpu2NgC1tbIDcu9O1tAUUZwZ+fHwCkOKRofl/iVGZ1N0Ld8Ei5hc3vI/ey8Ny5/LBIZd/1KUy9tq
oirIsgf2tAy8NzlJpD35jFk2jZaL+6lfA19IF7N+DIMXp4VkOseNIDS8Z74IMnXrPZWQiTiK5PXJ
ujZllDriNvaXxlHDCsMczMc4VQM3wdEFRAoOnI3hSnABw4hVCZReWtjGJ9vKymaeNYzoyHeddxGm
14NyCDZNIOwlP0h1UJ6EHgEOkZmk2Pa3iTe69sjrOi/qAwqTnd4x7iFauCM+n7BRQG4ElncCoibJ
0vYWfykZdiubD2pFuAVjeCisjHytDDb/kA3DLokFM+AVi5WXq2xCIGCC4M7RdwfoYKUAZLsYWhFW
7mzr94MNlpURq+HyskTvV2Q1vdK9HbdwEWP1+JQROYeHhkM7MjBnbl5gG8JEcm6ZGgUA6a9KpNCB
fkSMDL0vYutyVFpUQBloO4vZiXje/QdX9lmtUVIU86Ud9dC3d2D8AVi378prWrMjs6qmsJ54bsMW
VfaFU5eAa5yYNzYT8g1QRZ8dmZJkp1V6zcgFld7RTnDSYBtcDniqlNJWAlIwJKWG5GowAnWNULTZ
Ycw1XLFvRynTUkLGAE/KRjzoS9iTlB9xUpD8EL3cnbOYtgHZxHN+NmD6TNoZGToNU69NkBzYh/eK
uFPBtkbqxm8FblqIAFWFHpvFiIUupiUeCmqba4mA3CxPUXIRX6fCvaZhr5yVp3qAJbaZWkJfpBO9
XvGtysTbYdE3BUH8JYuQPl3Se5LjDKU2jRNRf1wVl7uiP0Ytv2apIvdNzIZrde2sEnL0olSXDKAc
XWNoe6jFPbHi+t24qTD8xPRuQwOC8/eJfzggs4VQo8YkDBgXmxnxIx+Cw8LXBBffVOubj5XmzJWS
/Rx9sK8aMDP/0+Jby5TecYLQvPIIo2eo6K5ft9fMMPT0Sij5NbEVKSb4TV1Xslpvez2r4YZvp/z3
2y/C6xWuT5X4EyRELSmi8FxRu0IRTrbReyPUMLBj+PU+jm4N5XehtxAH19hynFtTXji9Iy1CnDVp
YyJts3GkEkb4+Nxrgn4QED+3lHfY0Be9mGIinMWfFzluYkpNwylR+5XPSjtrZJuK8ZUY6x3tUrkS
zFEbgmitCE8O4Dre0VF0N2dyUqksGNN5kMXZjgjWdD0XDV7c3gZAcIniobzRFvQEntW3fHqE6gTJ
iHaAcTk9voZOawVy7Z1S3/nXhQ4tnRYn3UNgVyLf0qU1JuomkqEvdk91LKW72ndEhUlnyI+Vz/YU
QMJXxwGkGKDvQkyHWJlf+77LsoZ+D5OK+itktxEYmwQDp8rnjTfYvC3TsPw21E3BbOt5z2YqIZGW
c+iYknaT1RdO6tycjfDVhWoIgkgSlFrAcKDmx9DoSUCoJuQlPFTB74yGgFOyQ91r9sdW1U49N0lk
p1xujYyeMI8Ao7/S6hTZMsiuNioXRUXoFAewANpB8qn9w7z18s9GhGIOxhTCBKPmS/gfsVzSXzXg
e1lqTlm3qaZIYiBmR89b7znwTAekdpDICfH+Dec891uFz7Zhd15YG4PY9xdegWjKHveUAaRzng4i
5JDx5GPihG1MU28L5ql+o/33R4wfcanu4HTAWpQrbR76CS/NWzWtbNZ6CkpUu0alKFUc3kMoFz61
b/cpuHuOXz037X/i1ZrAkTk+y1asZ8SPYxUM58gmEwx9EvimtrRaQsew/qsvUq12ofWo3wiCAEjV
ckDX6XrW073s0T67AffGj38H64NrfP7/ReElYE3wMLqKlGcbilQrncwb4pQgX+QPDDp/1B1dbo3V
GQGvQFM7ctiyRIb4AdXQ/OC7cgrpMpUGdYZD8QWcQ303gcv2D6gBq3N6qT+UiIL7UXp56llA0Z6J
EM8zQZ/24wYgSmM5BBMIgIL44orK7we80pM+DJZaNf58dIanXA5k4Hnhlyjl0C2sgSa7WiJcY9BH
F27pK2Kf3Oy0NmESvvg9v7tcYOEz9xcPjqf5+t5s1bTW1MUDWjZYTu2HA85fcnwAUprOCqJyVhTK
rfZWwyL8h/RNl5LGiss+p43Wfc568QsFjOHqborGsz5rkTAtEq4z+K7P+1US+0qFDwuZ8u/q4Qqg
buoZcxU8VAfdlsLxxxoA9Lb8K795FjhOr7O76oFmKuHwXbpge7BbvfmIXz+WkOS23HYPLefHYZnc
69Vps46axQlKrh03T0gJ16bMLBRa/2MxxrTZ59KLXGKpQOHZgEBRrKQdzZ1X1pugh9ZRLYMpSbpA
LDMo9tj2oWXmQ/MZeWV/an4dUDH8byHvDn1iRL3cObrRV8VudO3gPslzDJJIb+guhNLjf2Qug1dT
yh0ZPmft/GtlGSPcPt4UiJxSicYo/Dnd/IHd/qlaXXg8PUQAeQdrinTz7oMfCnKSeGOgjWm0/bjF
mUY4CBzaVW1lYUJY1Y+GnBjeiKY8HvfuDKQxDlkKCjRKw8iKtWOKb+4hJoQsOK90xslZd13PHr07
BpkB/T6ZQ3WrxsowK0uLxQ4yx6j/PkiWPQtvd9a52Mnb0J71s9pVn7ezPMJtG1lWZ6VxF2X4TNb1
s66s2i68M/u+actUkoDJtjUeAZSWH089YnEcKTTMVmnWLz+dPoYXyAEI3L00Ae6qTXb4PIDwRGPN
vqPXMWwPjBh5nCbC/7AfT2WdwisJFBlcVaJfBsPIIRnW9qQ94pR4FGKu62gH1dqzP7/CBTvm/C6Q
jR/PDv5s74p5IUp+wdhzLfmpVJpgUUP52oFC0mcLtcDJaZy9ryvz8Qkt7bswROsURHCKYmeUO5WM
RdhZdIr7d5EPSwYGeq7QHksvWERrYVzA0sebPqkRuG+MudcRlW8eRpS9ZinySnOo4a9hOv3BZGX4
LvoRto1bGckkyiHiN1m77Sw+kDj1sefqS6BnCJ6vdb19Ssn00CX2rZOpfGxcasyO04Nj/Ilnk4uV
O0m2FvEfAvfUgL2MhJCXFNS8rEhPBjl7dDxHxW0svY3NgLJ5VYFY+1u1NSLjWWVBPqQEREVZN7TD
mbBNEXjxI4fm27R9MBiJg+mLgv8fCVCICxsSTddDLIqKpk2rYoWubJPJRANQdDbKdj3G7bgHie6b
NUWis1YcxVevdsCKiPnG0K3hrswzNWoXR7H5D/FsHct4HSfzJvtiBwxcQoKzoOir5CfvMsI7Yti1
qmdpNP7OCwQHdpeb4hJOkN//IczENnu/oa6QgDW93rSn0+ITrU7ev8VuZj+utwHTWrov7gkFbZJ6
T1KoqNkgGX9zSQGLolLxv0ldnt6HIUV7mkWTayg9jHgR4qDNrhp6skCo1tBXXhFdNGO2JGTWxhmH
KkrLU4tZmzS77YVPNb6CkVIo/bHXlsqRjX8QYT8hC4eWUYuR5kiJ47P2MLXSxIZwuzfAxL76pGCv
i4rMaKtzvfTSHI6aUECLr6JPjAWbH6DjZRPqV4xQgrlgik9oi+uxkg4Ux0DZe139efPpsJuAdbMR
I+XQvHYcVkGDz0TId0usK0hOK/etJxi3yCkX5vZJoiNpg/Gvw9Y/ololm2S5ZE25bjivXT6u8sas
+rZ6fy1CEoMWu73u596+WHIyid4Yn+fo4MHM5b+cGOXV+mkAVWbuYyJm7uhP10V5tgdghmc0CalH
v/ROlrjPHuy338oByIcNu6amJP8vK0zevWyWdihBorP/HHQGd3GNoLj2C0Bd2ZI6bMWbFzwJ7Ffq
L8S11UdQKMjpT9SS/iMucm3ZKH+J3RoLORhZ8JGglng3ObHdDff5hOWsdhCe27Zo9xZem6oBgrXQ
Y7QJoAkyij7sE57j9NBO/XnvjfqezRNa8jvEKvp9G6DxsmzEuMOvR9V7/U3C8Qb4Zuade85ddHSQ
6BZNz/90pABsv8MQSPV4HrmaSbF4aZne8buANrMxGg7M0u5QoToMAGGLjaOy3/csWD9W4mlexkct
HTcMkZZQgRF1wjHXcSl4IW0nNVmd6mEm39XTDw09S+37fUUppxTNlE/0qg8t1FOLqv+CO82obbo5
GMY0C74hqHOGMDFbrXR2qsCXaJgnwST1IYUiHj9Xgf06mUlx4yeBhZR1fXBN5eGoKEkIgJ9T3n3Y
CeYcFYlS+gI9kfH7rxA7WM37l+gLCQNNamm/n7R5SKg0uDxEXRypAXVsHkqVstoaMvm3AI37qcaK
s+zM/qOvlLlOidal2uY667GMVrz/7s3JscZNgCdu7AY0Bnv2ok2r2B5X26vGOZI+ogpoBewZYxKr
GviOViaWxqjXU0Bh0VMgwuOzh6Zc8r7Ih7a77krCo80rzjLlvfjbA4axxfmK2Qk/AlpQHg0NpsAZ
6IYs2UjTp3nYntLBcBom3TQX0rp5Bm/tc1pvgdVsUay2SoFRQxYglcyBd+gemXIpIqFO5RIR7YZP
hwiShL25kiZLZKQz2inXWGSv8tP4gqbNTusxUeav1IuDADhRYrkCInf9kvO5ra9jaD+lNLl4QY2Z
3VIs1xYgYwgK2O+UHtxCCcdeRcir55DS0EBiwZXtnRtbWSZ08ZICauV6YI/mai+F8/qNzzUqAPab
XzTE3ClL1TsWaZB8OBIwJ59cbfSyAnn+nJtrzmqmaJxMZ5GEqXCp8l9B1PdkyPZVxkFpkX/wmLWW
f6elqAo0iZEDhRCYvGSsXvrZOotYquU7A8a/vD0A6h91uhrOcDyMcYdHtJIwLaDAKHUM0g5RinUd
4RdwHkAWlaCqEJSTIMBJUJNHnFSq+Pi6ovQzSdqygWGExPKvDGlYBbLe86tEGIqQYxcLFa09BqRP
VZ5uvPVLhLRzNBbce5jGc+Bkb4Uky/M8EuGZQNxwSlYeeaGKKywcVLBnDwt6YO86fM/DAqsREAYa
MO/Q6ikOltwHxjnxsY9voMJ+uSshtPrqA+Mr1+h0O3AZTisWcXxyp+qwoYweslAzLuDSPqL1KXRw
6fkSw9piV6ZqHIqI3gr1nuMSix+mnbpFZUeOg0NnOkZ14/LSY7qbFhHNzaV3w5T2iJYvOIPzOFdh
f1QlHgWfroipvRL9lpBk9yPNmuYuqC33VfaYx0BexAvJKKe4OzfDXrH8Ce5NCXVWY7jVOmKIE24f
3pu1ShTW1WxtaYdtSEgMYtffKEqRyTXiamV1auX6j5kSHjal/1pzXZWAbYQe1F4foBNO59/lddon
vqv8LTl3NnBmFB+odI2nXPz81h8d1dROoH4NFqqdONog3X8GPxaDeWBV418lzzyfO8nn2T/IMfLt
rrEa3TcKYV0YyDqEa701xeQnT9CtQ78dmErfcNU77X2vE30lsD9PWvrV87YaMoHUDOiSYLC3xE1u
mVlsALOaS2uXfrfTNuzWUPl8DaHTDlot8kPHz7tsid1zFJ8s90G9gdg/FCZIVbdMgx3nrI30tcu+
DtUzRPf/FguVT1ahSFcbfMbAQRGukaN66XdEiL8h6s+i19imJLDbm4RNrM3p0Js4sEnNsHe9KMPL
4XRnMaxoYEwH7STj5aSlFUdZjIEph3e+SyRiKV/je/1AsgKT0y8w5h4SVlvPo8oUtYmTVphxR2AB
H33szJ0zZb22gUvomi/cw9xAVk22x5gQfHa8KHE/gbg+zA0egsaf+iTyDzgnkjAESJ+uUthpWIr7
LFr1RMb84k8PlNy+Zr47bBtLLUqsRtpMIVs0a7HmvsFYYNBqXaGSxgbL5+0Sx5ufxme1P93cFtHw
SK8s+ZskfWn+nqiYgXmTM5vB8GXBNtY+KSz6wVfvqKz41Eoo2nPNAnumhn6SFr8FCbvBWwNFs9GZ
opzYLNW2KSacFj0r/UsNoXhC4CT9L9NG4ir+8gwoZBNVVeA17d8CD4fHsZuGp/azHAIY35Tpt2jU
oaPc8MKrrFHHboVaiJmGQZDnYGjRvcQuUZqG0X7jnmd+Q4iQkPuLK+GJiKJnoMnhd6sDYF0ApWri
mZ2WTaF2bWRsHRQ1aHPGIGfVo1e0bSYCnEZDCEY8eS1CLk/iVV1c1vYBBjFZwyOYyCH+lHvypiXc
OrxiEQclpcBIhQ44u8NoysIsoThqVPyjvbx8hPXH4xmf1vZGhFRk1hmYfsgqM0y2dEvxmNnpIATx
TctrlC6QqpA8e3BXTgkiAAGWBrg2d4MEcaMNuVb3oO1fkaShlFcJjM4NxCP9Ga7uNnKme93cx5eJ
GTKtIJWb77iuJhEgyfjlwWwiImtYtWTnr1fcxBXkY7Y/J1/nR+XjGcLboJ7g62I+HBlfjehQ9rWe
2ybkWagb+HYsl2APTnOLum8TMereAe18/fX7d/4uPQwOhaagOx9DIx+7a6GUQjzvt+ZIkNV5mg0B
+vpiwhuEx5sWjEtBOCHPneEQnFBWi4noz3eDQAFRRcEl3AXsIxnlq7tEwNZayzUOJ7MBCijbu+gL
0uqQKGpxVX/66PMXFjaZzKCmI5dfq1dNVqqHmgVlCYhBwwaBvg5QzZLQf0osFA91jYwH78XmZmtC
GpoMZwCJGFG2mgzb1HbW4m4vKrM5yeCINZCkYpuBNK/6Gy1xFxdTriLNB1FtrkvOoap1Qayan6Dv
XAfa1oKRods34EBxeT0WXY6R9hsETr1475kVbam+uOrxDAzefgHelF679m/7r7Jsk1NF3ATWHr41
FqicCn5qvm4HBLy90WjpZr2IWEt78p/rUxZJEkM2YQ9Vp5izOvK+L99M/33bKWBiP8hl3B9ez0EO
h1K1cDGnYjhEDATGk2Ipw+u6CmSLrac4pn8xinZ5hwctGA/AGTyFYSIycDdKDRa/17IUyYiVAC44
7Xz7bdyznpMwJPxmubIz6IZ5DKb+YdjduY/Vb7brQshkeaHh0ubkQYnvkjLJP14HyTGBFHyliY5I
ZXxbwh9i0nHOlvfy4C4pHNTrp/N3zTBMbaE8AQIza7g0sNVo/wxiDXGpwbyWIqwcZ5zLUPCrV/jb
cydMMlmgLbFQCg2QuLdYkBKkEuyBaF2NSawjspbohUAQQbep0nHSnbk0nCL6viwUPzkCnMm/W3EZ
URC7284RnzOo8PekxSl8sZzAODN1WIJ/oVarCz3tBeRF5bkR30UAMQerUYBuw371vBZT9XGIQxX+
HXe3vssjpGHl5LxQRiMury2lvg9Fvd9unVd9mS6WyEpJXZyEpwI5x6EF/wnruzQ7iCruKnrcpV/1
3GAY0Kzg7jNGuzAmo5whcEibl7SR1qnFnPTqXsuoIe8GxJC4k2FMitueg2QFCe76VOqSo1rt+2mF
jpEWOm9vXOxbAjARheP7ki4ddNrMOji1b8Eo2dePM09AN3ZN/Fc2/SkQTrfZcqYiLxZ1f8kGrsh4
gc8JW26IwGsXO6j3zLfvjWRHnnhHCz+avl+pkuaCaawuvGpY/t+f8sURjqi2ecofykI9ipR594G4
uScgZ8bz3bH2xmO/dYF7omMS77hlczsvwx2E+E/j/CckmmE7VKYwFy0P4wxpDEP5GtoMOwZL78s7
cYCOigp/kZtTkXmhCHCL2l8sB5HBmyXtDaXeFE/v3Q/M/5Hr+qQP7PbaKp/1EkLgSD/k0KVIlLRr
XKdgAaOUYvkyeRpgHEOutCZQCXOVwP2mtKlVWIvuuktmpqBOg0GZ4YEauUYsJKJttQ/PJMxzqs7t
Ff1HPMJ1L9FBVrkpzeEjgSDRRjfDZX9wamZ6pfElBQ9Raalnc7Iosam//+e8kvSOxd8HDRg/gTQh
u3E9HqkyosLxiIduBcnvQnLuoohyD826bb9iRmQgPBdhxZ2Xht47o6+fOSARuzOjV6NItTbLkxSg
LBafr6UYSBhR7zD9sBH9niChJiGzQSDYH5tZO34Rfq30F2RIEpkWTCh47TTQQkTJfQfTu0kize87
xMOG2S5q0//Pm/a8fxOaWraKVJeaCgzy9XLYJJL2CdE0DFNJ3Xp+xSTr6XkNOttE/PM3LquNATvQ
5Nh9Zf0UvoZGceY9LSsLgOfc405UAiIX+2MRs+3PusTKIjkqyAA401LPr7HyJ77CPP1JaBRCX97N
T6QZr/EyoQ48v69CQ8m0eWkFseTMKcJL2x9qLU8rQtvc9+bu2x753E4OXwiLP7Q2PDp60kueaaP0
9VJcR0Od22NJCcmj/zrgYAhZ3raPLmD8RF1HhfX75ddL03Yc/6DuKwaDRXfIcpttHcbXfftBQVRY
Syo2Wqk1IITN2BPWRQ+LAhlZD8Jplw1yewFWJz6gTRTAjAl2hBs8tNIW+FwoRjTNHJ/6D47uJT0D
5GozpxRXYd9dtpSdKLdctiOsPQIUP6u1MnzuGFFCNaXBuRBoPSv8fGSrbDPdd5wqmrEOlsrChpup
z0I4P64eZZ1EhG8n+4Z639pgSJo59iHES32gOOWEf4CvwRQpfgsRXv2c6cRPx3fyqd8+fOhVipK0
EqqpQ0ewtd2E9a18tDZjQ00G+8mtACZxmlKipbPxgsoQtchitmxzrnkyQ0o61j9h9edgqmxGmzje
hjgN/XLa+80FJuQV2culMlJSBqtWybs0Y2O7WO1O1PK+fZgB/IfvtBx2ZMkrWShdAbgj0TYmEVBS
QOpczvcY9OAgW1irZA6COV6ytVo6t5OdFuQS53crpX0cwgHD/qHDZP5vhg89yp/R5uQIek8li+JS
XXcA3Y4u9WcBURw178HamKRDb/8Ra1LxEV9pABwBcN9LNUiORHU7R7m9GKkhTqD2n3kSg9atbjqL
CYMxW9o+bQNJvEuwBTZPsLzKWMjOGDaDYrwSKVaUgU/kC+TZxtkQtb8qZwrkTKCQj76NvQEQy9Yk
2NVCc6jjiWpWAkr+YZ5/fHe/aeaHHKxKhE4Yk+wdd3ZLzLwxRnD1EU32eeURr7vWP1fR69sfwdyD
7EsUEVMfLA1T888OI10TkXwqlfWtzKGrwUNH3klWFIIYR4MWzVzf6/tVW/wb3Vuhk9YoCHH4M5oU
8OmtLMoxafF4YKqi/26GjPqNH9xU6WrBxMbgdl3CiSqv6qkZYZwlbuAsU//u9w2NNFPTfIgZb0o6
54Wn3AtuY65yVHNgLO/ZcJEgQWDWys09Q/9a0FeoB+5m1Q8uLe8HS9srrm4S/yfuRLAD87B3v/5o
r46aWVtZ7LYUizSXvEG/tms8O+ZvzRSYFQGQJIhVkJOmRx6slToGU1VcM/Gi4ZEke+8XVpsqyIkZ
Vw6UxwvI29RDdeEyac2n5tXAwCSYoCR6uJnUgkMWbpvZRH8/R7gpzOlB9k2QJzuBOPxPzYK44O8z
LFeh2HZjJWnmYtiFvQZQXMKMgvddzi1x7hBOO9E+W7akJXq6Ayn1swdaxpvi5Ehacn2m8jb/dUGm
qjFhmCsspljFOIYMAtjhuoihgmmbd2SCT/IS08OX9AGobGMFmSOxE2IZ9pSYw/hvE0WK40TlVGJT
KnBQy4BZSPiBALrggA/0TTe8EY89mi9JDl/fqreV+Blh0h7RBPNleno/SDca0ic1ES78jndqlGyB
7F6ZcHX3ZVDHyBjzIIXaBVkGaVdQPjr1p9nTQ/+q4K6scwQ09vtIc3OkfulWmCQxm32wb0Qt9VfJ
zGRYrKnferYYZT4LTo+aHX8kJ1jx9NE7o8i/mQ6/4x6KUqAcRsJS6scXh9fpbW5PagRtLLlx7O1t
ZRe0vb09E0TC02MQi/zTWfCq811YOmw0e3OXYsnrcrmJOm9Nrm2PlW0kFq/h2NLMJo3ZQBot4aaM
8TlplsFv8BwsLKIshWoTXK+6ynjooMbtSyAeSDXlP0yRAtsvuxtVlPc2UsV/qInDFpeMPstswXkn
h2vUGKmzhl9DrNCEv86SW5w9NnMgXM2s+3NVoIWHkbVZD51ojN+xd8IeKhW/0oULQ7CD4YXwoBNF
GsSVULQCtzBqc5IGCOghuJyzbblb2dwW+O/Y3Xx1pU8pJk2ZFlwNyUfR89EJviert/QNYPVQZGZt
7rPwfZID6J/qew7/CdykY9spfu4mQS77zpSd0Vb4gjGe3NmUDuL6qAPMuxIZbbCIqRh+1Xu0/YGr
waWNAQ0ve4QEi3QuIATVqyeWcFFLwV3579aK5fK7nGXum7hUUkrVe3EyXgvlx28/sja+FlZxIEcl
+E2LobFc4FAk8uXbpZSqnstSpIZOj53ZMbLdjhCTOFAdAcTQLgnkQ5cFVNErRJJJtvryO5ZhPwPQ
YCnYVQtDXhBj+rsi+MaEg00kBeSBrL0tJnUyltBQrSxHK5FMc+JSZw0FEFKG1XNSG1/bWW0Kr+RD
CLoEL1qjszlteZODgwhxPeIg++wWHqnZ9D9Jyb3SA1DHEdNMwBb3addeAZfMNxqF9tKrVAijUcyH
Mxbu9uTUa88jX/F8lK5pFDTHz765U4GA8k3dTPnYi9gVSlO08xpW/Gdqlt4tRlWuqhFEqFHP9wtd
UhHsIIAGuhP6IEZTfND/9gw5lUwA6hu+YVSlHD0mOFfJryV0VLpNb4ziRnSJXJVA3jptaaCUALlk
TGV7TOAaJUDjEGruR/qy6NhcwDNOpJCCdBK0ov6Ag9nGzTY+Fb7a9EZsplUWz/iJSpCjS7wSj0bl
eIW7z2TBJ5zFU9NJzyAtiwbI4Pse6FYX2P/1xH0uDIncsRT9g0lzXV9vUIy2MOoIUVYGw5KfyBAq
YNFGmPOZj3ajxaalf3qr4XSUTjsZurvAO9xgZTfVpoHWo8G6tEltUzokS3a4zEBtVtDy1oTRIQG/
wnXwFbW0VzIKuT5rEAXwG+LEgAj2BZolSe604MAdFeXTnLh9BwIXU7ruHvdMcGbmL9hLfMAZqUUb
Uv9wsitHjixwDzOxmzFYcnGyha4j6QA3Dn1nFqqffpLz40tLt75MsjqwmzI0s7MyWN5/GCa8zrgV
YLmEvifGoEd6WdJJ2XGZ8zBMnqK1ydXEzXI5fDWeeZ1nS0xopVPkfabVG1LLgRI+4FwscE6GACc8
B9le0EwKqP5KZ903d5oho6CXqX1s456Dv7S/K9pMNS3dU42GVfRLwXJxmlW6VLB4MSLVl44USQ1H
+uFztY1590bB1Px+N/Asl2Md2WqpjsuRRb08Gq98jH+w/cs4PMm6/HC8nbQUBtiOF9GNFGXKsV+e
DOcYBTDB6Kb9rDZ5UtL7FART/aNY6JK9phsXrEMYUuUDVsFmJheu6niiQQj8nrcHAfJNqanikSd8
b0PbkQseq7XTH87zYhoARg40DVBQehIE2BhXZIawOoAMLJEWpKW5gXxTJ85cS1PHI1VWzzd37q5V
HLcEx3PPjLw4n42SN5JZsE5ytK99yZ8B0sm40k4xXJz3zJxh3coPvZlCUbpaQPpgEiNoIeNc1oAX
d3XInmPapCrRw+qUs570MTq41l6E+5zu+XOwM/YEjsnX4/QuTkKw7hYoQyLofI5r+N7Oz88oWzZJ
QTtJIaw1wmggsxDj8PVJWYXHN/9/O21O8WI00gYv7cm32fifXzP6HTNltrWXMUTrtAxoonQ+GQ6U
1tHxn7rnieSYxcXYUVp8MkIqC2Cr/8Kv8S1ksR/VXwlnRPHSTv8QzZSdGeTUxvdNfnuTnNB5Ix78
RBMVaOtlg0efbHFHChxftbSvr0yaGGgOpb5S4Uua/d/Kn9fIJfEBHEpVOM5QPQ3E7VMaxXRbbmLn
fr4VjniIEvfvHiTYQ1YuEVxCCA5O0H1GzkA10dSJWXexn+CvGAHPaFnm1ySqpR9ijQa9M258KRoK
8/MQo1YZ/RuOqPwN1rqqrwH+AoNABRZeH1QNy0vVDLpp/uzJbiWhWN7m7jkUdO+W5v0IO08i0GT2
nmFiKpI6Eu4gFuzKJHCX9JyCufV6SgdkHTgIClYfLVn4NiUAlbZOj+TuBI+ffjg+IVyFa0hM5Pdg
6Y2+HRat61zGEOVFTnvSDF3pybRJBun1v8k9enKaRrwBQDNDw//P2EFEnhjMgsPVCy7Rh7kQAkNi
PgC1DQ0gJTjYZnxZCvUXauB/+/Ocwm6PPVc1OOFnh7OEFeRAMtiKBMvROtxUYwBg054hMF4v7rL8
avSXr+r/tUYRrO/NDjaQPbbSFT1kmmbWT6EIlma9pjnQGi83+lzUkn5u5OgW73AYi+1mPt1SONwx
hSkXR8Dj9WE38L9eQQtFmhir7Bl94e/tr16MYNbFXUjh23dq+T+TcaxijVbVuvixLTUkRwCAaT1H
pRIL8RmOf8ZxXxEANsii1Ubthbv/HZA9o6LEVgIhjYZU8+Pq7aLPWNBeHmD848xMYdMA4m+epFA2
FUiCmsORBN5bTNtPSLXKkw/XErVq8yiXkAA7TU0U8LkwDvX/G5LqN2rYkK9ux2UtgPW4HFW/Ldv5
InqlcBVxmvQgjNUN5u18y+Igz6/qwsV0O/V+Mz8TiHtBfiLzOiF62bDo70X4ubIoARBgWrDdPtTU
/VkoqXYwR2JDMFFa/9jm+u/wKYp4BgjCUFeCUtroprEY1qC7b6jeZ2jhPxi2/MKlzl7MjV/b0NPx
2B2y59uIApSsqq1X02DkaMGNqLKzsxF1qnhj5k1Eai+FfGbyH8A+12JF6yERs+aHJMvEV2mzCwm2
70kkb3HGTtaFCEe+WiJ4xdjHfjjFbxynHKQP6SNZdufD9OdM5nZEmGP9k98BW4O+X9BTKV/kKWfI
o78ePtr42iYuhSA2RuG7S7WNAgGXPXQDczdtJcWwb+xjVhv+E4OWRaCu7eBPEkXahVb4ACsoPHz0
8F1y9tux3uB1Bat3KbxvQNtNkuZdkWdfu3q2kdqkYpOTWxjWuKxSNTx0hSehl2WIDSRgT52XZRad
amPE5QRed3Uf6FtZUPQE4kKP/FLuxnaw5RvhqlbTBWjUtKYXsLHllOXnJvcYuZz/h0jWm8b/3Pe0
gIBtGIYfIfCAIrwPCzQ63ogu60IhiCFt7JTizWUpzRaAqz4adn7AI3tDUHuAMd5bYga52Ua+A7E7
oLWd4bASL7Jz4papUGK55N5F5TtxAv5nevT5uNiCbLS9VEoV5uefns2x+52e3iueo9X7RYJ17j/T
5cbPG7T74PIOc1ciIX72H6+ExIzxFt7xJ3yJo1tDeOEO9Ur599fvkXB+geDba+G3aoqZMS5VmtP4
Ckj4AqOEyVraUENhxEr+L9l0LfBuD/nDkHckO2gwX3eHhvQe+8fRJYCVZNG7a4/E1rLSUvIwGwI5
WcT1UyGS53Dptfvsw7PB7pWR0c9bl6xakG+YsRbiPRmD8OV+S2VnMwBU3AZR1ip+VpU35BHDVbNy
lFrzFngpMSjQlAR0By/JvJ36qIbmNJIDan5qJp0KHS6fLj6mrcW0SN8MjuQABdz2gkIgTuatsI47
tx5ep7e19/WzHnYZSrXLm6hXhDUrXyythkIwxJCGJ/hnaCPpdK5vciJkg1DAw/in1JSvfnDHaqTX
B83JRgjmtmuJJ3C9l3MYQcdpleIc53inYIqJ5+NcN7d6VqQCVyJygBmL9Ri1XQ91RQYo7vU6QADt
oGkZKpPA8dr1aGM8B3rhl7S7Y1ZGvQT+CMF5FzNvtTTr796bVmf6sGB/sATM/4ADdbdBnV7qeEjC
hnMJxjB4PodHwxoFhe+jeKipgbVzIUwp0E/qP82o8TJ13Ofmdmesvn6q6uTz7dSyWLvuOAqkZXGw
lTXtFMv/87ur0kL1xKgZ+fGu5kI2uBCmlG1/SvKWzI/tfOaXtHEGmQ2zAJP4UVmJL58NHMFPKh6K
LaPD3rNr1D3JePbAkewwLbYJUw0e5OvdnSzeNHHnY13ZckQ0Wpa54ySiY81XAXoGn0PKkqtke2ra
xz3zLewIgNx8rz+tI0X4nbG8jszMaTr+vW2sbkvryU5PfhqV6uCVt1GYX40jdgY/gMACWKaPldhJ
VpnQ96VEnc5y/zR0muSAkImDLog9qUWE820mlIhE96esq/xsykOVxnM6cahm2RqCvAA9BTX8g9If
6t5SBXBch/LgA5/P+mbrQU2hERK15QTOtjaFAOgU39xK9daKG4JyhzQyC8XGjJF0FxofK0fQHO20
9iG6lba09jr+t+LWa9kpBWJb2MFOf8ina7BT9EFGPaqlA1Z2iH/daDu0RtWxIIpUV2WzARSLFdJs
eQjGyYJQMuqADpp0/Gc/uhz3Um4F3npjcCBTFe1Ke45KlX87Lk54J4+BoUGyBQOK8QoHgMAfIDuD
tR73OOlEBmxrFUVQ8Rw2Yd/VHQncA5tr30J9J2IzVLMahmmlcPFg+WvCTYkpJF8W8UKmJCJmrjqP
TSZTSZWpbicVbj9kbH/Uew3P6agfqTU6pQwxPoDFt55AGRqMU1t5VpdiJfUKrL4Sh/xRJdYwD09y
/bOk1/ERBjEIqNXsALjm89VExs8kxUHfxCMHDPFSP5HI+u03rCJ5AGrS4IfDEzR1F88IXUJUDvjc
mwEWGykSSN/1wZ7xi+U8HBgqfQsO17ZNtxwQHNsig7xtvC00seP8gYWtVP+aTqX5Notpq/Jbg/cZ
57m2c+HQ+QYISyY6jw/J6ywCONgW+sziUir7yTDwC7N+Udt8IsGcDse4jOZ/87MLiJGk7cyS/4Wf
/Nm+HKc6nqtCQuRDnUtfH0jSMjZYvCi7Veh/kEkhFXJIymBXUPJ6EqC0r3H7jspFE3WZs4qglyPn
Zrl7QyjHk8JimftYQKAZ4p96NqnNvKKjdhf7yfmTKIuv3lGvSnG3crJmuPiW8g+Ji25rCE7qgKqi
7bPh1UNUwNczpcELg4YG3cLU16eAPgzwtCGUrGeuy0ZTAdoB9MsWSju+xLM/VPeosNJZ2YnYJD3P
ZfnqWhVYChB1eHQDqZnPNCEe02nSMoSh0nfZysfME8HD68pQRikYyZmZP1DtSDxqU3XHN7XJmhnG
27aKA/2mnkr7VwQmruZXCzYepzzuyTIs1lHiPD2hmVjG4BRwPRNBBlQ7/w05E6qNSY/2Z/OOAe3+
cpYpPieEGuSwK9p8QbvC6RIW5ylRbhdh5GhRHMmfmEiTHLP/0dj7GzPSGHFMw/tcNMUJibl1c7Vh
vEK3qwHgm6LLecmvVZYjXcarfUOl5+lCfFZCKCRSqUj7lqTyzdgLBfHbdXaFYxjqLMZLnCvLBz5Q
gchcHDT7R8VaSUNj9gElx4jW6x+Gf0XijE+M23Dh90tDMAh2JZhU7t/YzbvuTHSCS4dxWUFOPPme
1Llq3nZN9XBsYz7AwUhYJQHE57fClsiNCTVVH+RobmM1bFo7887FshNcHUDBo1m+6vWS6AHg6PlH
9aabsSW1YglIHC0HtdfFRjmwCkOGWDCJbrahc/e1acE5BrCbUSiigg4RRmH6UCiiu1z7d/rfnxYU
fMzMo35qkMlVWRT8zJodh4mDsLWViHArunqFZ32v2Vx4M6yfgeTDyl2Zn9156TCj7n0VyAfYviXj
jgdvv9+YnB2q9TuIn4sgYzdwHaFaujsmp7ILmqTHxUHXiIZ0Ior3l/VK5LBLKNsoMsJooew2C1ND
J+SwlrqHFIL1J1nzLvFfIvqlqXu3nB5lTt/zfCwsO2UvAfVWSZJRocp0UZoKnfJjHVRd3BcfLvxo
EMjuGN/afgrdqzhltMC2VQT19rJaM3y8jVFoyBzXlbcIEgXk6ltMabM3yDe5zfrU6bmDTEc69dKu
QsbKzaccG6FvwXqkYEvX1verxwXkxWoD1pq3GGpoW72Ouj7el+vrAO8AUlXmFL1S5Nef4vqFqwFm
b9++EU5+kv6da5aQmtJymnnJMzP/Yuxl/Jyk+ZwIv2YLJmgsqj5sgPlVYLZZ3x3D2HybXxxTB+gz
A8i6wgsGfxForklnaoatLqH7EG4cfFg2WQ0y7Ehr8XpL3VbvYArWs81YJI02y3rV1nim9VjExNTa
PAn+SCT/Vdy7xqe23l+Fd8dKblGcmct5mF6Z3tYwik8hHDR8hdn+ql4cBM8DnT6/dZpEBnEON9kK
6b3yN+88adSGqzeku9qe+5Nge8du8+mBR00/piwcvhK89iqSfKz00zDilHgEtQR69vfAXuEshX4Q
n4n7Wvx7N/3yYyXbZPoEvvt1yBwTOJhLp6jAbV+rx2+GklIsTHMftROVq0yBUs/W+ZMjRGB5/0UQ
fcHE5gY4Iv2oCLfng9Tyzly3GwsDUxCj/FV8xQaYX87ck3FCLaWY51vhHlt4So7+e8a5UMSAA6b7
FhRxo1obzAOr8Vdvh0485SheaVetiK+qmQbkEGyZVNJjKFl0vAfsksBz61K7IyBugiWbinJNELjg
b/rv7FZaNqAOiRM32HeWsieiy9Mpd/8iauHIEnPBPeQ5kLCGzpiXfy4mIHLrq3m7bAe6qeoLfg3/
X4kKe/SW4oRIobyZT2XByRsh3tG2NbXgNGE7bkPLCKNKAt7Elf2C3hkOyIQo0/YqZy2+PyN/r8AN
DaDDWohcU+sHnGqNYJSfTWLaGPSIJ4FFeLRqQiXTHQZjKpLzyxxisZ57bSq11fVhJFxZhuN9NH+C
fO6PGhYqhQb27XRYHRh5SGl9BhHPkt+F9unkjpdUG9a6J6/twkk1Op2vqP/2IWJrK5wHBXVA6Kc+
JlRg8YUOQsXJXQTEDtNMCP/F6hxzafsTinPyvsB6+KSxxE2f0lnERKKSec6LiTJHJ2SfgljxG3jO
UOvbFEx/unPB+1odFPpAkqEMP64kwhMWUT7B6q4DalguubfrA9s0SprJuQVD+HxNXq6TsEew8MvY
Yvv//KzNCIpqJf0DKP4dFJm/e/XAlpNKxnIjzY9z0vEnqRSzyx5MA0gb+3GMAeBTxJqhGDjsPgF6
4foBvCnabsFcksq7fJ+qDaJEJl8FXEbarTXS+RYxR4X45M5PmSOiRwGNl2vJ/McGcp3bjOXKJVRr
kiYuea4aiK7QA2kHtURGdXUWKqECwRVmCJyajZM6A0jwmTBZ9VM1CVBg1fkQKSi3qNAdiDrb5HA4
99sAWddIH6I2D+cAMdwyqxcKEZJF0tWYTWkFvP+rsmkdLqAYyRCUgX9oNgNC/zHtudqVFVvPL2FN
jaBJL+WS7/JqpSBreIOmmlvty+yn8Lvx5+zSVbjDiLZYc0aRxUyOyf+S6zTZHMWMSa8LM9Dmt9bV
VIzlvx4by+1M3wLJ1Pd2gRh4pHz7cqMsmiM4+eR2Gp5NhP4xFQYHgmUJMZR6Ks3XtcSGjHCheOmh
TsCkz9t4S0uBg0lxng6Ad7ei8YGq3gF6IEW+gCrQ+x92S4PcC5Ow9r/TvXGGYwfYrvUtyj3uxVqA
TsqfAE0QpVtUkHEuG6cvkt9SDxclNtEwDgWB6ZThpJjj/9NhLbg81rMAbeoCQFJJPKo9T7PPxWe/
Kkrw6uNZv3E7WWXbpEk0KjxTT1oW8dffp8zYh3IiuaHj8smEt8Qd4JyPTz5ZwYljsspTHs9C3XkK
4Aa0nFvQ0o0HUSXINCbQTuUwzd+ws1dzvoX9VsitNT1xheRM2FbntWA8CcjGQdrIHLzfIQWfeClE
SAhsULHizHsDY/pCpztvtAsBauFm4mlbq0b/InzTgt6R/l21stYxuc3RqSYj+mfmp44j+TKTH6xV
pfMEH7mtekgtw0N4euaOcVJWxjbxxjyCCJK19vr0uz+PgDB8xwYZUJcQg8Jnmh64VxBsRJSvZt8l
XfoxZWKxpr0MCnQBto6QyKxD/D+N6DEM4iMNM1fo96VoUOb51jXDD7XES7QosCPo8VdTZkBjw3LS
cgFmFbNH6+QnHehGcKudao6PMhe9plyDkx2+6l9HXjiaVbqBDxNk39xYgSQVPdkVL3apc/DJZWQY
T4Bd/j4jc/OsQ3IapEbhQsPMLC2luqLYHzjKuHiwX3LT/RC6yyhz/bv9rqhX2blR5VEmSmPx7r6d
xUhJEIuBtDgtbEDy+uBlyNG7mItl5W51/ww1Zm+1svUPAGNJUc0mWnKVVNOg8tZX5M/+D8J8gISA
wnzTEza8XtD96AIdvVAHH0QU8Xs1k/3W6ScnWAhx9Z3UWQaCt4VFVcQKoj6bRV7lc0mW63ap1cLs
AzIjRMM7aQARdaplOiDI7xh8Ag/546Cyb+gY33kSKhwkt60eRZb5CZuDB//zfnmkUf6uYkoE1NHA
r5X4+fHNHtwu26YYIPFUydbBm8208fLC7vaQKIhoQRv8VCJHPieNKuZhDpMKrmXw2v3nBL7dx3Yu
VqiKbrV97OTg1hN6slyJvEt05Z7ytnCU9AWpf7YjxfSdV0hTj+bAn5Di/R83yOsyBPBI4lhIPo5E
PxBnm0/+V1xB3YBGa8AOw71X7WowmeGoJ3BiSlWZKjnztwzlunA73KN1l3B6wgZ4JHci7ftRKSRk
uvEU9F2/lyhkHn57RRYGMJbXcV2RwzF8Jlo25q9wd5eIL3GNE4rM+SFJMJv8Co5RSvd9ztM8YRRh
GeffgCkBJWxfahWwuXarTMQgyl2+DdN82cMO7PKEPwAC/9RB8lLAUZ9T3gJgAPI3TwRFstdOl8/h
e0kmlWyMFNbAYMo4WciKb+S/Y9jygJbCdHscDL/rt8wOZUooMkv/9i3KCs3pfWSg57AXuE/TMUoQ
6B+cENAllDyX1f+Ljk2cKc+u+0UNkMjwWD1XO8x6m5bR6p4rFytv72oKIAgFFvKmT8XyycBnUogy
jrEyLgh+FPvVtMqQ16lHUJfJobF+LKDm6OQXFCab0/T6R9IMaPnLYniYIR8EKnEYebc6liqT1EE+
q1XMlheo90IH98M4ud5xJDEFgMTMBTdzrZEIQdrVNfroAgBwsGrz6513GJWTN4T013yZMRu24llI
EWQI/Ql0X7+AAgAgFmiXPqF5Ye77JssexUonsSM03NtoLHnstR2hB7HnQIbIOhz/Z8W3VgRbjbnd
jKTD3AATsKV7xbMmNE7r8suKmjNvZsu2GRJ+ppDH++AfMEH52lfurs1ohWfjn3S1UD1PoIS0JcYP
sUxmpfmekZaZ/D3LNGQPAcuHw1sqIW+OhiTsrhwsTLIInMg8W/Y+dD+7gqPwAiLB69OjBkTrt4PO
GncRuZ2nKDiEcmyTKpPhW365ghdGJSEpkFQUg7wwAuWfPOKDJ6WoOfysnLyuJFV4rT73neGVZP4Y
3Uh1klD4cZubykbQo7MfD/3l9bSATAOPZ7dEx/GCr89I26gexxgtzVA8463JdCuP1RN4QbI4Hm+q
OHtiUEw6mR81uA6oKwJzEr2q9l/lMCcLBCaQwA3bsAbNf8WD/8jk/AhZnbyydnS+UW7wJwVACsat
dTLRlBGWUeulHH3sFcD3rNiabmAgJ8NTfdKPkeP1JDcxxTUFOSjdQ3OYz3vJ9msFxIz6y1c0ftO8
7whvOMmYzOJVbiQPFi3SWQnDU05nS1EINml0ko46IBckMUofvhdJVFMOJtcr6ZXKD0HJfPth0u+S
gOVx/n5DrVVE77BjXOjkNhoLuZ84En2M95mP8CkrzbfdFBiILbbz5WDcFK+XW7NLGXlABsh9/3hk
v5fvHIxQf52qhxL3VjvJksFy/x4sOTQOYi3vAo2shumlX/XUnS9YJv63rfnfX9lWdphaPbLVwbfK
HL7cyCw9M9vqvSYoUgTQFu8/BcQCG5Fo/sbqMrIrn3k5AGiTdpEDZJF3YDWVsrqb8G98Xh9gfndI
VtHVWDs/sSOkpIZwvuoEHyG9mZdMrUuw8/qTOIHp5N3RJOFwrIzFlSbp8SOfbkFfes4HHcJDSk5o
eGbgs09h6DYJsMBxO6lJrg6/olDx9YrDmTVUEOW02u2EHM7cnmd7rjo8HEzqfe7nsXs7eeQMAMxU
5BHHR9CiC/A3TMy5Gjxz8AmGCuBQotMoWN4jzPZL2yjyow5yZb03TK1of+VaTGiHWnIOSitov7x2
v+jv04gXYj0lu1Zkxy7P/kjUnNLzzDAj3Crou1bOmiQAWB4Tc/dzyMbuvnGCNGkVwjJcG8ePLe5Z
vysw5QApDfisRBTYw375iGUZrp5apIyAzUhVL9Ecg0fnW6vuxvkTWUAo9ORL5nctdwHHIQb0DiJv
7LV0Bx7JvhdI/Jex4a3xQVfz2z5fgK3AZ16/XAyo+GEQRnP18PLL6IcRpK0wbQngfB977H6XW9ip
8l/Ki3c86toKx0pc0qSg/4pgVseSQ6kY9egEYwL8Xt4sNYLdpY4+gQiNwBr8cf3X1va4mlqTfz6w
Q1BoafEuC44mmyYl/PQyxkGv3aeqBfMjFAgwSWZ21I4E1/dyFJa+mFei4ba8NWVrDAYzq5f++GCp
5hlKZ3sy5ZTJHfFE1UaOPzVvcIdUkOqMObznX6ZQnrLJtG1UaUpLpcELW0vPu3Z5NJOIuopRs5FN
c1mUR/AINclC2i4XTCboagQ05m2PLpgRrHOwWSwwDaJ1TTAkyLvxMw1MYUCa07a3nuQBQeHyk4P5
6xjt9DhwuvNBlanwZA0qnywBdJULwxP8hilcnl6Exlz9BkazBpJt2dr+lgt86zUIiYTDVan9dMKH
BAaoOefkDv/xzPZ5gl2ZOMOt81X9ntUHNCeoIPuicVExq46cfyADoK4ZdR4Ocb+xW2YXNDixkYqo
Ngdak1aKpOY9TQO/E24ppZvIS6V0FdkAC/tXzgRXZc69wMhkDqk+Tgpu5ZsQnKDd4fvJ6jM16r8l
JuPe8OB/TbflGPzKgU1UBVoFc51Ik8LeZprHbVkaRUOrHkM+nItyokez+FIwkirnv1lSp+Eg8iVQ
RE1ILDx1Fk/tcb1D7mLid7xRXTQo0J3OEz/U8JdrW7yNCEmAxTT2Va2q9aue8hWtUkchFAlY76iZ
acNxnqkqKBBNlcU0kE9KWFo9bBefMTGGXk/JF2HNSPQUqSwMWk3biu43crc2U11UElVPDirrufg/
dGCCK6mKZNQhj2TQ0QgYceyhFbBGrZeYuAPxAKGJU5eir80zHYHVYZTA1HjM/wAxj9ycYLqv5eEI
l2edC+ynk6/WnHseTVKOexA8I5q6AjkHVvJM1SqMGwJ9Vo2hbwfI5twtEdSiNSkzdvLnS6GoCkHb
4eQ3kaa/fsc6XeafJhVk3cOvBhPFW5vN4Awt2dfLE2eaoA0RVIAZAElauliWINFSM/Q/Vn9uOaK0
SA5aG7EhIyCi0Pt9F7SnqY3nPfPpHuCwLy/qMTFb+Z3Ps44NH6taMHCOvs0l3iskMe+1yQOSTrZ0
6kJ+95A7GgraesGWbE8k6pDjQhr4wmFp6X2wIA1rV23Q0Yw0SSGrmFqv68fBndwsA8V+1rfi1Be3
RW3LhPaqsxlYufkyYDGUFWRVPxYw36JsQdSXL1JqMW+mR3hxXQxJumqZCgpRDT7g1Cz2OKUpUZCw
rK+3WOabA8/UdzJv8STgu/KWltH25iyIncKUneaCPt1zyZCP5Mc7nJBFUmqi6eIWhB4SnoS5ww9v
BQLz0mmZslS22LBXMYjIKF9zW+1Q7rlKuuDWn/Xt/KA3HuumNm1fGXAWJ/kSr7O2gFeQwyThT00m
Rrdtt5RIKOgPDrQu0rvwN9GZo+Q3W/MnZD0lM7JzYgEGELwVnoE2FZes4Sbl+rr0h6HbgwAos1H0
ca6MoZgm7Sa7w/3ufi5rGts3RjP9225uT5UGcEOrGjMHjq0nXwKDxoxfFRyJ0KZA/ZZO1XmNZpz/
rNI2FPFJ5FcRGSn9rcldezFRxmcZxZxBV2MQoiD45GEbtH+WtN1EG1wdxlFHc9I5q4V+wuzawFtB
gNl1aQYZQU08Whse//158DEOsXk6z9hBq7oramOPUQVBdi0dZxUBqyXWG2UavcvBPvI+IpGJLiZ/
lx+vn8vPl6uNato0yCJo/DJiNs868a0j5jAV4UQeLMfWpmf1UnyuZQGsNMXC6CAEsnAChGbY7AQh
Yvz1LkdwBVhhaWLX5X6QxkF8p6Ji/gAdXOg+MpGArtBUsx7DT1/ZJhFhoW9NvnP7Htixk4j4R1BJ
1PzpWtVqklWucOvGVOJvPm7zDBqu7h99715GnTM9UWO4Rgf7yG3eNK8T7zLmu5XDHjCYEAAoBqSv
z0eIZEJ8VwUAy9TgdV9Ugyrspr+U7HBGTlgs/AekuuahzPWp0/uNLwtAxW7P5PGFrHhd0cyW8al8
WvHaFUd+AH/bNZW8b0Gu6eJ8AyjsY5EQ0ZYd9fgaMl1Opupd44DBFHR/RNGIlOWP0RnF+TZY1jrH
sa/L5YZKnlvks+sP4rcI7OXp9KCnIXOhrAhdA8fthK1ZKlj3A9kaiTDejtI1YkH2JyC1bWcmmtjN
bAAjNNfh/rUvEA9IW8UaTsdqgytaQBjicExF5Odu66K7H5k5ijwISNvH7gamG4w0wICjfZSzsQv+
+lQOpacZzt/nUJ7+JLIt6ny7QDIAjyuPv3fq5q9Y8DvOu6rivEXpDYT0427ofbdCI/X0j+Z/YjxI
NP9AUzrDTKmQ4BJupzrwkzJlJFemvw3AnKE/Kftx5vgNzTu33D+dp/4jIky37/KpeaOa6J07n6mp
h0DapGFxVwnPakHy0HoYr1ANovvoYSJ3D3D9xfr+NSXZ43rs0fbRh7kamoplaY2BZpOXqZ6V21ee
gfpevmoZxuv6hZJ2XtbPYS3MIO9v89In8XXGpqYMRItcbZQyeIk3Oc/f6BKCCgvAXYKjPqjPRA6w
W1bw9frDEvFr1cxggYe7gptyMB/dZLpVmL+PJaqRv0nrCgOQ++fufSl0C/0A+PRjWFqnbbVr6DMt
wYiCOR1KJ0xU7O30l3tbp/Kv6Y9pPH6ym8X1GZT55wKMMSE8xqLRrreb0K2NR7NDGWu4tSwpYC6j
K7jpmPHYOZMxBg7cItH6tE0SJ+cnPTKL7wduZrisMYzcFyJuBNUpDY9BEMIRCwdEqLdf5oe2Rf11
HJOrSlynxMle8AuTWER6sDg8m1z0f95PPpaL/mq5Xqv1t22u/9a0n//PzvG264yBYtzCTHDGuIho
NAcnwodC1sOUQ+VjvTCSePqpgdPcqCH5Jc+9Lh1MS4p1HoOcINvBUdsKqdN/qCJbUZDnPykOENdD
zSr8LMvVHP1WrLEiMp3LBcv/Ub4IBq3DycRNtFEh+MMXn8IJUW1jJHtFAUj+/kff2OzRY/LrB6u1
sKTvqWp4A9ADtWdxjFUXHOBHswOY7+7Q1xTBVzlgME6BetdRyWxeVIUwev54IbteKH114SluV7tT
mC6Js24fv+nKEjVeYQckzSq9Nd3cNanSKi3YE0MGl4QvOktYPUXqqBDei+ctWtLIzx0A71dDTSOC
prQdURw0v9Uf2yuq+IpfRao1wjCl6IdrbGT7c3do9M2ClcXP3h3Qkow6uv6Rkpdp4at3ntbpkP2x
rwDgXErV4iarXVWZ/iBFQY7MjLW05lJZjJCt4oTP2LF7A5eoDPaQ9Puag537bqd6jgWnLkl36yYx
QOHAc3G5W1CuewUatNy3xLDw7ItjIkMpu7wXV/haq4PDsUUe/iIy10MMPfO61kkSuK2lpr+CehFI
4toAm7jlmHJToqWCI2pWJ09onYuYXu9uOSseTXUYSlAPkItgvKup18MmwWiELWqeGNaV70FEjO3P
UkHREKc0gX9DYGoLdP0TC4BUqx9yXSUGfotu7cq4gDFAS1cu+tRQjcX7oCUMHdqBxHJwUXWgv0vy
30PyPSx/P4gpaR/oPDZT9ivkLv7w4KZkMNKSV3xgy5SFdBa1eSH2QzAVdUzjbX4NXiGcaDDwx97y
OD0Dp9L5eGQTcLE8hepm6qaIBT9gOIR5iAQpcdoq53lWZZkZRo4s+ZfeVHd1kqfcx4HNuEtxx+1Y
Mq9STvFfK3YfjX+MHLQvPU3itse7tNCm3Krxi5/MQeccpMzCUAKwkaDY1248E94rl1NPe4BEZkVf
2KIe9hs7rqMbfV423oUVJCVTGLS6h3dumJJbhgW6JxAui2uuWG07bPpCP62x7tFsMHahUaGBtS0e
pMM4YIYH3zZ2rvunZY/PppkB0/kmPSGtZuzC6ivPOGvXACn7zMJ3jqFudVM2CZYskJq7uIL/pnTS
wNVeXaOsAZoJzTnfdWtpJLhQhZgYONTRJFBt4qwpbEh2pVOk2lzbKgbhEZa4yd9kG2q+XwO78BXm
tAJpAkhxKYi5dR93BnpHdEBvoxx6UrpJEs3Glf/DgW7x510zTjWLRcxHfgm4YkSdyxNENRrYoDNz
M2HpAQC32nWSHnp/T/0XZj/sc+ilxf7qHucylU7+ztcvC9tNQ6eN+tXqWdX4wkzMrEuA38JoT80c
3ehi+vzvs69ttICPvaXjPWqEr4AL6HZM2aSFaZSeTvS19Q82hKBbkBT9/t0tkgaLLlIZOoFMKi+S
tpSSLLrcjha7lxBlriPe00L+cyIiefZi1/rQVZrpYXyyDYMLuADjXE63u6R46kSQbMNFBe4RrYFS
PjU6P/VD4/AoXSvEVmvKZa44v+5TAT6o7A5iZYOajItUbBX4ZE08pkdQlyX01HrW+VsKnuo9oQxa
Mmtpe7nVBKGauWkKdb3IhLmJqdIbvKLPoyalYm3RMsFrSQNRa5wa3GlxmZHH8P+sWfq0uozhwGXA
XlQodGC+SiCqWNggqI/y4IdKlg1v5pZEWNAvvadAQF0WuQkxb0hY/px0LX3NaLRVsUjFBLI5A1zh
cOQZOTZ/KiHz8Aaw5da6MQJutSyp3+HvHy6SNQif8o+lhnXMmhOmGN9LiCR+vR/1F9t9Kbpyo5wT
BTZ35ceFesq1Q0Y8IDbJjWPUzuh8gAvrTDBkWT6qquMaVQghoZhtOazmvQTR7SpFW08/cKZ1gdgk
FSynINcTM4RxEIAY/ryfRRisIYKTwOEpQTDjX7dqvGhVlEYaZd9hhf7KgH+mXC8VBTN0lzNwotzu
4KcdMeKfbXzRySjy91qKHmqwZ+ish/FIvVhp7vaGfm2JJCE2mL8YRRU3OQ+8H6vMb8Fc9+Z1h2/j
/OCD+h2dIyvQNLheVqoGBMW7LX/sMymqRFRo6sPHPiGSQumrmYLV+uGfPlkGF02RdGx91tHuUurM
pEbDmVeuhxniER5AEYCKbtFnfPTt5XrxjVMVRxULtkG+ZP8CIAgDH+BZ0PBu04NrULKifDM8Goig
Sc/LTKnbpfYHVIc8jjXT/JuWNMnhwgOtjg+Jsh7CtoQ6yax3brEWA6bClYK0UVsSxXJPOKajO7HO
4eyhoNxlRb2V2tK/z1D42oSv/KcvmIqc/AtBIZvTfFeqPI5kaSZwDUl8nNGrormhO26lo6RssQmC
l6ujGSANhvtu48554tUW1PcJqrMUYGj/i9KWQZ2GtbhzUAcKBBpS9BIx+tXViF9+CJFkeFGAf3Km
IN2fb2Bauf3zPsX8ECJm/PI9LzTHsxuSlU4+21J8WwxWu16VUyM5+OsHEeJQ3XAzccLkE96akc2W
pZvlSFjAmqokBOnZyv3eDt2Ft5oPsvVtmtoAn97Rgv/83+BcCuX6g6NbtO7zxh+b2PsxsM2Mn1uW
7qie+zYcFEGBvFyN59t6+8V+T7lFyIom87AvVXzONRLaMK4sgZlvdYp/yu26aRj+NQxTTPK/lycI
35ovi/PflAW82evKogGNl6aVkUVWlRml/VC6GLI2669/Behk9xhN5b04vLE0Spow9af3+pY4aSPT
WpTCKKMkxdbvjJ2JVNAD/wINdYA0Wojj7HTrBj9FHHZs8Us9nrEBj8t+9sZMCx6WbWfpddllfDzI
7vDORx5X5R4vVL+fuAMCuNEuzIZqGPnVDHUao06n8+43FIe9T60t0VyIvHyCaD1ahd8KhrSFzoAc
00eAyKw7bq8ELf45iC/EU/pR4YObI/Xyh3dh4sg2vjA/swXY509sIE0F7Ha1Ut6MiIr3YxxL7wvG
fmzefe7P2YPlc8DJwMpN99WgUHeXo94TdVveBzO0x/HvZMtay39RMadYwi25o7/lMTaatsYLvjg5
Nr+//9n65qz1vwPeKjXFBS4f+H742iP22UYUSEuF71wPudLo1mXCI1oop+TgPqmU75p9ll55xrw9
bD5M+nYU0tXNonpNxydt0p5VRgsWa2D/J4O144sJG0qMuJCwm8pwuhaTNH5/IN797oRkcMTNxfvg
mYd789IwqacXPZgOqJXavc0UYTaZOMz9WAA3TBL3H5P7dyV4Aq5Nxb88Vk9nUQfxuTOrff5wKZQk
2JPHwDUjS2hfo27ZtimLIMQ1dhw249UpJTsSiSMrzNYBgT/WHNSmlsZ9bHfOzTSQq2AZJfTct7sB
UCEu7kM+npDoHP9LLzoTrunlg2A85gNf31xI+HlRbO4gpX6uDlCTMG3ILziYlS2oCpMsmwU7gSIC
l9fRcUoabTcF6luSELfh9yjDuTIV0g2v9tfsy2VKu8tDxKOr6J/P7ibNbOrNWfmfviWAO35zrHap
gVoeeJyIazbz6AepKbwFO8JvWAP/ZY05IKKuLZOa2XZgk7iGfd/4C+OtR9S9K3LqImtWY+a8Wskz
kJkHjqKMFPSkcc0W7XSjOy8J7kSDezQ6li8oWCt+pP2YztzYiCcHaRzjNLNnRrFTlW76tj0aD8xr
fVBqMlCd3BNCIwfAT2kXB/crqefdUmG/5Au22lzjsTj9sARmoF6Q3p5LVKrWoyPWJMB+MY2wKibX
++RSne28M9HTbd4NZGNIZOwthCMhabz9Ix4vo6jTlaqvr+I0GSvZm/dyP+Ih+vflO9FrV3LATSAf
f2rd9MscIfYI6Xojll8f9xZ7FgevNwZw0+txcNsmJRbbgpkKLceskku6DnDBoPB7E67sc7zD29He
n4Q4GtKBPJc6I2A55xkUajaB2LEGkojIHJHWGo4EZMEfIftCmDmiWPrRr9YTbDkgFRjgc16jp8Ov
XKWNhrGbmQJJqBGTeLOB6UKhOFpGyCxxAsOaSc3jWWtSaRsX7iFbFSzTtYpKRZcp9LkFa1iEm0Pn
1FZA6jU4euxr8KgNJQVB9xBbfMFbJNlNqpMrT6nsNrvfktPqTL4GqZLWpmDqVvJhnXAt4ZB8/r6r
cLH1bbC3tGxplbnhUwg+BYmk/+A1FfzhACFbTn0+rLJJ2YzPdtXsc/IHNUX8iRTuJYeYTe9PYg9S
+ylbgOqifHWfojLjIyfHfYSuWP2OsBteR9M71Z4r9uuM7Mu+5/prEb5duAFRSIxsE61jQiu4odGc
GUJ1UI3OXF1FCNKlyPfeQx+IAnZpEZhSHMRqier1NdE5HropG28JOxJ5A7AQUqVAlNoLBkto9JMn
1CjtF5DJD8A/JBMT2YchtGkQT5+xNUqg7HrbNLOHUjkqNvuL3Sxx6Bw2WLtt9G9LN2m+m7vviJHN
aRE2WrDWoZA7iYpV7x+XhnYKbPepfU3Bp1YfnJgn9NP+ItkQYS5Pe8ciKTo5KNndCzfQhkjm/CWR
jAeltjiFkhO6puxGmOEhlEs+ncqrrRozfgq7QVWYQ/my37l0pVcIg/qWiVCtLzMSMv5fZnL+XWqR
YVVl1Wt9UuelMBUZQbkTFnUhbRCUuZzbJwBbfy3gtGJEeY9TvntthPfXlsdP5v/GABys2+4tdEST
LmtMrAKk/O6HoYbxCjefb2dKA1dSyN2FGkdYopFbo0y+kxMluU8XljgkELTm0K1LvqZa0FasDcTk
SpoWOXvhMtaFj6TdKCCFxPtq/cOcvcUFJxn6K60cAwaeDh6S513Laig0ZEl5yYDqUhjbbtG7cEuN
ZAuV1lMNVq5DPA44ldOqQ9JzfqrQ6kBwAEP0Sc84KAu01/BZjlxY8Kt6tU4bkISJB7i/Ql0e6jFZ
hCm3IK36Ml+aEP3M1YWzWDtCooMSvXFHAm+AAdeWE2BetxgVwoOGjTPHfCAWrrJniri1w2+7Wn6Z
O1kvWy4yTFwqRC1NQYEDgQf6cd0aqjs0hn3t5TrmkdKt5bn0t5VagfdS8XKFboVflkjmVURQ9g91
tLC4cp3/aifZTef9lZptioRa4XC3n6lnLLgNvQoFpcAMuWAAfJYbSDui88Ct4VPMVPwnViQZApaH
uVzEWG5NkBqt+BLOzkzYh3WnhqwWoIQpqpqFeIwZqIoJf/hKYu4O0ZFi2PltY+oITQn94q5VdJKV
sEPjKoMjt03pR83QjheSBxXTaQnqFARQFDtIqrOIXhn+7EdQXdI8jNRAyv+yiUF9wihzm+p+7ids
nDGYcgAcjLtGXCO3G6GxClMXy/tNILdGvhg7PLs5H3nAKIOxF9ar7k9V/JEHAVJPQ3S1aM5hgs5n
6xWGTCJVgHAo5mw/x2e+MdRYG4gi/fRoytgnp/TpR5sH5Rxw+zroqjaED5ReS3oHc+vOuAAM9zHw
poiWhCIrXKQ6tUFF7ZTiAuzkRJHaZ8Pa/kfNUfqSTx6+Q9cDsBvV3u0kVkVcgkGTCrTFx7JutlXu
L/98lfTmxR5/aR7Mg64lLzhpljh+bQf5foVSJtFJmLJsJbq0cBnMBdcIjtJJYwsuouMQUwYPbLkW
STHxW0zt9gmrRe4O9HYEPd2ny2a7cWkH4hzzjJYf1mPzlm4X2fHWpinWItaUUdu9HZWUK3mPD9la
vt19dtrEI44v2tS+scXp68RIv8I6sv5i708d3CpQwX7PLGS3zKYLXA7MNzbpAeGHMEtdsTaSC/tc
FoGPwH9S3QXCyatVEQhxG38KrxBoIv38JQa4oixmOMpomzRfRSPBJtJ2MEkqjbtimO/oHDVw78Z2
rGZAe+tTIjjhkOfpFnzNksA+FKs8stMyYLz9it7VrUyVtT75Sb3WZNUI1++4pjWSzWaTEeATowx0
8fLCirXXme9tv/a0nd5WJoHoN3KXTAZ3Is2Aw0V0o0JohB/4wQq3X693iCmTUKGFinUmIoax/cSW
1WDl7TsxwCM9TGXYG9OwOBkQXSb8Paq/xGgfdWx/8MztETP68VlTmtvqrmn+2wgPUik1WTWN1b5g
ArGkeMcUu034zkEiz+zsQgj/NKhjv50k4l+0UcbV3+8tgFdXmhYWkjO6gXopENvbd6N79ReIiF0w
Ldu4MuVtLyqaaKxhhiUoD+DuU0uhIH5YUQbGgrmPB1PpoLQez/RjKp+JGVYIqq9brtDn8CU8JHqM
GmIl2P4QA8L8pjJ8YPUoNDNIyVbT6E1PYqGHrFrN0/i8AbSBnQNZHSUU4Vaja0yZTwNdE5Cm8YkU
BCI5GZOkJCRd56N0JrhrCCUr0XSpSYrW5c4r7xHLQsgciMXDXABZs9qzkuexez9erGzVcqZjqAIg
ebK2izso9eGQK0DoYmL0TyJAFVXuZGBbAUUUXO9fH0xNTLS+R+HUC5N8T7ht8khNLl2eMpltqb5x
F65nJuPTBRU0sx6MZldID1v9uQznXHGbSinrrPFUX1850TvqfB5h6VEW7EVSnLZJooQkXr+G68PI
cmU/IYLFdqXohEqU/FfUo9nkUmhzFTDEYC43yX9iipgGBc+nzWY0JJcENaI44l/hPhLjVOzbA1GB
qZHx8j1L45I3vUyJfoAuffTXkoUSYLDp6sSw+0T8SgKeJWDFGCEBXu4XbOKMkfa5aKkAD352Avm7
MV66Wtb5aAJmmEd9cjjwAzde126XT/zyLLEQECwy8Sc9bhZSn6yXsUsNicECP+hkRCOKz5AQ09nb
eVKOZZF6x6brTDlu7edAHw/abpS5m5O6H7y0h25IEJVzBrTtGnjXnKc5McDrkawtcQpkONEO3Ots
CqoNSXtVYcG28m6j8SMI5tc3oqAysQjkBMXdORJX64YHF2e+hO43b7ds5N9l7+gTZMUItvxJJaOk
TNAhjEYc3+OtdjIUsJq+Vm0i6cZHlCFT5NprRVIbgINo2PvSGXb6005Sc/PHFXphPhS2SoYUziE3
uwei6b+ujs4x3c4eN6zb16YPVM8yzaPBwsLHZg6OgxNEENe0gLCTSYYPdY6/M41UAWBJ6TqsQ4VZ
V8eXSRu1cUSoryDVjYY0sHtsYq3h3R4MQe5eC3vXWIZUIHJujGsyzBC7DleVT3Ts0XtOn/ENqMiB
MkzxN/0r2S0KhubQtnBwpz4N8M9flPSQG5KQSJTj7yj0WOBppUlbGR3r8giHALBA/sOU2Cl2nQ2R
NgFIVn8loKanWCGBuUgMu5kqA+Z+BjxSJldYo6cFYAzbUc6v4qQZrZ7OAJyGIlbcSyw7MGt2UcNM
6Xmd0VKi6tiP4aklF3ywPabEn7iLKB5OBB+GjcwI6tZz3yYB58ox7T5ony+Z1C0256VHU4JJQdw8
YkLiF59/6pCMMy6BowuOe0HeQkfq+9h/AXDYl9xe4GCSBbmCjoeLsHbNYH1/Z2GfKt9QPM/GpJBt
SOa+lu07hhzkip6UJUtVIn/jb9lWE+irDhltVOkeQgcnYt+NUxt4WB5PaoqhogSxPhm8pWlK04Qz
6kA1naPTlzeOCX+G9SqobnI2cWnc53hOzrh58oPKLzoVH0S9b17TgPfs4Usg4tuOZIf5ARRufobW
wfQfT0i80jt9QaICpOLK0Kf1ftPGGEjGlr9PmCvLv26D4xKqsO7VzS34+yIAwB8U6+EyxLris2xY
RTN7vkOghqVmSaFDqpCaksVlEGSvw6QR7mCgQjbRp+Xq2LcANgvyCuvNNAfaX6YbT07ao7+QnBKE
b4CjdI6EJm8eX3Jo+LLGPPbqGegEvNuom0tG5xksFw8K5H+AaqJ2AxQnZxoM5aMzBgfUn6LG8sep
89a/CAHmIWuXuH+La1idMJQjucuTNiKJ8PsvWqMPN35qmuyPsMxkjJ+Sn30HGYbFRPEbekjmsag8
di/g2ce2Q9sUA4W36McH3A4yg6vlie99Xcv5fAmdUrN+kVta+zpfR4BkVFXyoD4Hw1A7l2Ek/9Jm
U/TkXjuMlSt6MFtMyy4m+VbYC3Bbg2pl97WdI+a/hBHwC+flPv3CSDMSXPFpVn+Duh0PLKlD0aRC
KzzzM5CvftIfHjF3VQltDEKoyhCOWmNlPRlNROimmlTA0EP/SYyv4w7BufAE0tg7nE7luNOn5fQZ
yiBwpAJv3f0kjVEUWjtEim7Kb5E0X0M/++UfB3oWXXFrWfvHVBYaI226u0FqrpjRT/7iVL5Rkd/k
Kt6rjR5DGkDO36a1rHzqfu986nY6AxQ9Q4362j3I0HMkCiO4B2X298ZiZ0zuCqwmWb3cIUQhq6fG
7jijKLQ7GtQ/3LlzBWdDlZVVgHeBreR4qWDrRU5D01iPMtnTH6ZrfG8M/9TZA0juyx7WvaayEKMK
oVdz6Kd+vPnehlJ0sQMkFnBvRDxLBSaT32+6zvg0dtXKth+uzZb8CgMVOHc8JrtYJ2ic6Ybg0jlv
VSGQkW+bWhpvjnRzpogDxeQxXd9QxODfjmn1snPBCFvr4jIZbWAdzUXSJkN/NJ7bqrM8dfwGsaTq
UmqjROABG0plUwHXevg6uNbChKaH4ZrDeA/HIi8Ii0Qj9CDcRi2SqPZAhXo3BK1NC0Bwhfw7N1Dr
YVaMYdLFiGO92DsWUEuYGHXAXHChpWXo/Ek9Jc4GCBuuUaUeOYz9VTDGpfv8oAsJddts2caW8mOd
rRpPaLJJHQsT3WN++LLWQTYh64JYorNa3CX5FawCFAjK9ajme7yt4ItuJHdykyQaBbsTnUo9cAzr
VtEhcog0JdLxreBY/JC3Sdi4R4ZeK0oYm00c3Q45mnh7qfVI1stI7Gyu5woXwDYy/FeRCS2g0BJs
TPF2Rw6SLs/dAxNPSnSre1SuqPwP0LYH66VCxE1AAQTZNYaqUq4u90No1xeIYGSp6zr9eZmum2Dc
g4VEfnGPBNu3JQQrKxQyAP888cZtWplXQMRO83oGRyDmQDI+TIFEc4N1ONJk2X5WRo85jNM4Xfks
MuvSYflQOMQfh8Nh6zXxG0XofEUVLZQ9j2P31lp+86YMhsVEM13r5BHbTniACdNfPYVdxtXGlsjg
s0j8uZaTibkn9FDuEWsQxS0dwwEPIWKy14OQqPMm1AspBUtlams3qfzxfmmKu5yVTrnEHhWxt8z6
e85KhMbgrToPrZBn7boFwD/k5pvdYQNXqL36KzrguCKxkpk3CFo8Cgo1UuZd0c2WSzK1Pqxh/Beu
3Syr6VtBwradDNxyHQVtdi1qAtyaY+QJb4ovHLVTlb/wckYls9OAvW01+ZIMil/RFjxyTOkjXO4x
fhkzRsOogyJ9/XtZPR3LNQy3k7xbuNe7FnyPoSctg3iIkbSVE09+2FCj/VzAdIGeUtwwT6d3Ie+G
ebdO10qzENKDhKb/mTpmCW94ih/M9GQUY8CA+ypfwjbC/rbc+Z5dV71MJ105QLqn4PBWRyWfsQxc
Fnj10cn9/iVTZ4VLRMkigGzUAZ9gtPjbzlux0zIThaFaq/l2TS0qDO6n6+TaGJ/Fda2S+rhWWAoV
wYVAM5UfYjlfuYIwi0Rsttv8itCLhqFYjgKMDpMNswzeEcTCwyCsg10ZQHNPwD/qDDZMgnGRZP3x
7kVbtdvIEli9qKg2FimssTStAltDU7P4qjyeqY3txQzaeV9SU423hPlsEJbX/5q1ll0i22eckjbJ
5GkCFJC3i7OGvqSXCLgE/ePFicxU/ov2mfOoqtdX2zyOjP7g2svQKZSDvdYvUJCWc2V5kuNyO/gn
Ldkhvjhkje3xPIa9ck+3qoRqv6ZDiAuH9kLxcqr+HeujAU43CxOP0ci9gMlTTuzlpyXX6Fk2iI9d
ITwSE9AhKjtTjikQWr1EOFrj3xP9Hyiv7/0+5kasAXEF4rlws7zIwVUNjBYcIaMDz07OyOXQ+Mm3
6HCKg/PDUlIUyp2hpRuJPLxnNLdxb7nXb5Vc/WPqYM4n2od7TRZthlkQyG8mu/XqGv8cvMTaFypc
yeDq4hpi0bEpavfktRu8Z+ewFC3zsicz+1y5bGb6Il4s2cX0A8sVsYfqy3Jz42U6BPbBWe194wzq
EGxm5AV6zRd32aY47Gjt2PVfNAwvNo8tmQ9gXs+9iFNlUaa1S2hGn3CTzWFKpJA28C68ZBB7n/UQ
DSi3Kb4eETXZCN/bKlT9f5atO/OlW9nL8YzygFpwP0X7F+SkK9Tw9pTqU9k7U/Xl+04mbDpu2Z0B
f+jh6wFsSWRcvonllZjKtHXyAkgi7Zsk6MVTQpEnTzxcQ3beVkjczRlZ8mBl+mtCRgQa1Z1ghxa+
3aYJJVceNqDJS+b2KnUtr6qwaZ6/cnPyGQPVYO86Fu6/tLjNKMtz03TzGOPz+4zumC5XLueLMWJS
+/QKMw291YJxr/hTFlOWQIcjDVlU1/IQjjd+N56bvkRzqdr1Yv5Lt3j0HGxms63IdVeRDQLlgboC
AoN0fTG5fWkl392oa7Vuj5Oyz120toCr0iuyIcRDG/CDKX4Tn54U2JtslEYI/fK7+TKuf+3BQ/Jy
XVz+U18NAzsbU+ouOMh62ohFJRdKkoQMuqCXUPkGP0U2ytt0CH0Q8ORRxpJHpAyaYqr/GrRTmsYa
SAejLs4Tr0Kn1XPaAbVyzIpI5vp1AzQJPiPzxGMxxktanx0Cr2CmVQWMtyks7C+iFAQIzn+oxNjN
YOzpRoR/qKmTjSYfUho2mf4ADc4C6LZcwgTR2BZDGH8ShOctKEBh6qmSr4AdsfBySO3wVyLKkuyH
rr4Jy859tfGJgdVJfCZLs8Qe9gpWaGmKrOtoqyn10+J+D3d3WlqtctODdVswmKM5jnk9t0pG/zMw
hCrO5rIluJKHkh1VN6DFC8jXbkV2wkn9n6dbDwJ1cdG8S4KyH5zOqgRxSA9jXyH7I3bif+yfrylR
JbjxoMZV00hqWPlxOSnOZ8LOq8GUDlnPeEip/zIDnOCbYKVR4tYFFJz1AKXZamnG4Sg/lgbe29ia
n6ofwtUVM/1B3kCzw/GUxvRQbaNRbUAsdNJ48VfzrvWnAAqafSO6QQ12ZwOVEsZfO4kPiPUKIc4D
eZ52zR6yMwxNegsT3e14mDlN3/PXFjUp+EMkWgVdJwYLG2TCwqYyyALPdlzQ03pUhMHosBqURuri
8juSMYSggcMrNydGzCRJB1CMF2v1JFKyJhp2RnYfiTJbntDuMO1x5MAzzS0hUkCwK/dT1gDMdSqQ
twY+UWb+CgfjLoyyG1RPwhqQzAin/SMNG5Xp1eLgPUFo0ZA7W7tiuRf7SGFGneowo1UOxMvUrAfp
JGXli9W4tt/WTp5L7LeeCf/R5hdMGwg4yBy9HIt7HorSx+VQ6Vfx6zI8t3Iz09KRzCw7EvXPVTng
EI+LI5V4ZRfCIYHdS+r8Z5YEhpvQwpPW+/5nq4I56hhJjw6cSr4k81560rSKadinNZtP1MmM/gZk
MI6lhw+w5TVL8LO5frRVowpZ+wefm13K1NFv5Bjeo227SDR23gPF4lrPXDx0phb/HLs35Nahrd5E
OFQqT6EwQ2jSrw1JkXAczmf7W0QV8uXNGIE/IATnfWLh9aFvsSgL35ydRtJK+UP0oxxaQIAgv8s2
UKUmf88dDMcrr7LJyqWkVue5iWKTZq4VBWq4rL3nasFEAys7TPV3v8llDZ6FlPtP3g6EhobUtg4V
cXH7YcKO1dDqbqgCZTLWnMLEyR8dhz6ahsirmPkhbBe+W+K5rZwPKKTFibZj636bVH7UsNs026MS
djuw/ROphHKy3nH6PE/DrLuMuDpO9tFyB0In8freF/aBsWR1Q18DJ3lzngvxD4/QOFlgFKm8pjAs
KMRJtwq8uzrFdMArarkG0Isj4lPsCZxVUoEwg0aaxlO7upALMkLb9NGespx1ZQiwzB+v0Ul3c+6/
MnOdnQhCwO+6aSmMq9W7w4XSXaUCOZNm64t0yW7zdyXPhB/rLyPz99RupkFuaEH9H3p997EEi1AE
/hmt2I5HfH8Q2X+1UALb1Dx/q+NIDHHX/T6LIjunN2PYTJ0g7U0sw7FYI0xU4ke0uUL1vBT4/8df
FiM9D9OQ34u7XJyMvMlEFSbtoemT43hNR9y9VX9hLdsMv4TPWejeIOabRpPAPOwsWbNRliMP0lHC
EnPnEViSODmjFcoceT1HTjx7xaY1AfemOw2R6U5aVjDxmYgqZnHrCTbPJsnbfCk0OK+PP8xBTFxs
2khipTqVOPakksPEgydUIYCaPEhp+VJiCYWkwlFC0pUhAkwpNI+O+FIKS7HwVkE1Neziiaa/6JtR
e9kWKfgDjBSLoj3rRdrG16vDGiq/DIL4YNXCRVgjJJ1VCixDfBuy9CVX7ynhOv9IIK/PlfK75kzB
eS0jlCDyGv1aIv5Nz6o6R1+yYHs7StxtwVewtQRVbOcXJKwf/JzwJ0vg59GWCGH/cgxowXK6lqLC
J1YMT3XhHUr08daJ1K+vpMSdtUuEQ5NRsjD/GMNpE6ITrzmumExuFZVgdqFvZDJ9WE7H0+9xzoo6
fWXesVf6pfUP6RvnDMZP4Tu454/b/LDx4l7eie9wwqMFFINC9aADKnIupS57PSFBZ2Bxx3lCl7+w
kO94vnUHFEgzXwHS6WaGRRNIT48yVT27JnHttV/OT2IoMdcPjpn15/lix9+kn1GRjkRnv/3Lr6Z1
lW9EUyxbsT9EGoT1zRR4oUNUWCg9stATj9gv/B++vh40qnLTKZ2h7uCN+T3Kpor1ySp3VbrCVRCd
Ki5IrXd0gvPUDb8awoVNM6htGxFjcJqKjVucasPBWRHAkCSH8IxHJFalBUFLCOemzuGXUAW8HOne
BPFUCAWdp/do1KWYMhbK7rMFDAhxLrTC5bvD7h6neucbfCVgxaWbFpsD+E5wZw1H0IlF+Jkm5/qA
k9ujA5JN3matAl2DEupDmXo+0dvxbEaR0NShn9kFbowZsAvheuvZ0KN8KZuc5frqwNRKxVmpZSR0
c9Sj+ThI0BC0FlEHYT5joahn8WlvchDFcKxWKPj9G79RTSI0Pso6JATzc22hjr0kX5cKwBRGgIpA
aCBUs/sY72O7di74YufhNq3L+jRFq3Ww60+Dc4x4p00cGl4M8sy4FHcX1X8b4LQt7NlzjyllYrDl
lR6AQQ51YV3GjN5ZJ2MeyOq+F6RNAv4sdC77nyfQvajdVvRdemP86dvZ/259eaqMOfMygx+XZvRQ
sbSqGTfhTMSG2OWi4SpK4ufQqgcT/6XU8aqzP4wz0GS89Kxj/GaEn7o5RZsD6Y9IEOUjx2MmDZZF
SBejbOklI4ukD6qkT0rUxPLoknUjzOiwERVP9kg78tmlvWcO5ZOSe5OcYxFWt3W6Svat4pfwL9G8
MEN0VlLqPZc3BBI3OfJ9BRgcENykUJtQYOySQ9pygXpv4q3NNK4HJ0//mSMtUAHtlNvh1NOLU/Pr
ETAREPO2KOok3cHpAo8tPvltwED9MPCSvl59RscNRyb9v38PddqzLaVnAjltLqcGiSyoDNsq11wY
3LqYXXex6WiZyuvqkBJM/p0YnkA4dbzUWmCplrCzyN9r7eCLEdxnEduZEH9eoaFDdKXa1aSuZ8sn
TzQQftBf2uT1lMpIpgOyfkahwenfPShUheyuzqEUXbaENiyIv42hY+oTKHUuUjoKNoMbjYz5GP8r
8r38d7q4+97xZg5QyYf2o77dX/trvHsIQ+gHhgbqO3GeE/JNynSXdsvIigAUiePlLgySWevdyA1m
AxIu6qKiiLab8q6EybTW9JPl51Dj/0mImwkMjjTcw9bmjjYyna+QlQbCbvNUiJS2hSZ8Gg6aUVS0
qn9mtbPC8wraqtxUZpy7tsvx3U+NsXiXKjGi2HHiGmQpb/rlUBgXARQwwt+KODJXn0Pc/2Il8RFw
Pakr+Q+D1MCsl3dF4Q7h2f9GyXrzW+jTtmIXN2P2gQy/chv7nEtIBB4UDfLyDq/WREnG4fzsFHnx
kb3i/mttJOukBLlmxEOgWlhPT/MDaCIz0OK8NScmeeq/ZhHvSJiOZZigbsEPRhB4YmTEsHG6lr8B
EqMleLCNDnUUifr5Ifv9GAkCk1NT0c0wX+dDlc/ivWtw0qo7xHoOBPEiWJn1fHywjY/2i8xmUdtF
H3pn+Bi1AUnIVVe6jpkogkDm5BOcrzUI4e0vFCIMhpktr7wg6oBFrsXfsfCYtD5z8nrxmR8bsY2P
l9/yrWjnTpLO1oUlRgrEw8OrclPo53bjF1ykUTDFGZz8cRvtH7IFyVdLoL4aO4/YXWjVjRtCnJ2F
jr3CWy8kYJ5vSVAGlcUBOwwHG3Wz54Jybq4FvMjNUh597+1OAFDmxq8brvOypyyZvFY5ebCCWoO7
sRBazETwRDq9Zy+cIwF6ehhy7agqbqpCsSZwVXOMAoTvRfUp0BK8FAqIMDeXeze9cTd/64ch1GLK
6ivX1Iqu931bCcf3ngF8AQMC4HI9xOM4i/s3grw1Pgzau1PbLZ7XkKMQyz5KZLagT4p9S8+lWFZh
z52yunSF68SZEzMemhLsPgRD8WuTho+oFG6FqhORjsCAeYl955t6qQeIoPvMDYhNeKN7xzCcmlcK
y0YyhK+koCltgM+veRuLLCNK6Dzc2rUYK9ot53uMA2VmHyGHPeQT3+jDO6+LViDCmPXqN2HGxqmw
BZ0PDOUN5DPuvVsSBqNZJDbIhVlyt6iKekXN5k1gJWYkj7cbn70sP1UaM6s2IL3GfV0nwOiKzn7k
piqMjeaRXo7T72bkHZk8Rqkv3/Bo1b5i4KF83zsUG5fqkBFzHNc9T7+d5SJmt/REShTjyFUt0SN2
+tj53BxtldlMzh2rVhnDn6SzwChZtF/DVkTK+/q+DCUgB1dns7jJ4sYBEEcJNxsta+j87ezgdZv8
5x2wp3AUvXvtPh+69J2iHrrC15RUIwdlbV2+xA8BarXmLDv1PeAlUmIFxwuYC9PSkaGgPFbRqDbr
haCaJdUOYxZWAcZF0awTZ6ZWvediluME0pMTUcvH7HKPkT/4IpCFavHzasQCIiw29dXRASvhnuly
HP0n4HbWd+3yATq1U2gMra33qA9GOVjClp53pBl7zFr6sYg3YdwtfBcO5iTKb5tm9lQklpLinc0x
xiUJB0WbRqRB9nnpKBzhJPTPJdinvcltJoiyr28K+b74JKK7RasBS8/KgXG5/uGHwbs30he1Bt8D
fg22KZ512c1e3HceLwqsTayAni2KJoBvc5it1jLP4dLk2oQyU9Fmib7mXm+QYgNQRPHsfbv4n+zx
GS+w4Mi1y480lzziU96ISVQxg7UHvsU+8ihmRhimcglHdgpSEgTAlpzS+usZ4bDvuEFGLVAVaMHM
0SjOUSjuVrtqqtnr9U3TEf04EZ5tHLTONiIjof95W1wcyzUH6kmIQM8DoP7s3ceu46XQ06Y5Rc/b
JPAinGd5muuiEfju9Ebj2y8ZCe7OGLD6sgT8TTkUrj8OE1VaqHkGVeWuwZAba9/YW2OO3rGnNVoq
tkv55wntmYUAg4qXtv/jz6wEq/mnE3LgOKhUrW6Xf720zWwA15cQd1d2xSGQy9LNayYRqx61ihpA
QxfXIz86+DZv3I5nZMjcX/xpV8+ncRltqjTuvknnuuby9C4qFoQzRgN+//+Sjg22DEjdjgBqoMye
zPeK9JMMCllYeJelREobeFJYyDx5Ugl6+D5fx5Dd9zGTfy3mZk1JcmU2v3vnUKa4ei+7hkGt9wlS
AFxwWdqrH5U0mCB3/i0tRygmlFSSrY5F5U7DIh1d7gv649U104B8yCUvQxbjwoz8Iogpl/T4GjuW
C7JqRKFEz4LWkqWmjgxccywhOhzl8KiPS/42fsvObvvkGNT8f6nGpRN6PbyD0vTbta6wYO/zCj5G
YJTxhL0ju4c2v0VzpTNf+LX1+CtV74FkFgOrvynsoXz5qu6haf2gFnJFu+JOcE0/DNIWQBl0Jxnx
2G53zd4VYDRpcyeNLNyqrdOeY6QJm+9iPaM841T3oGMA4OsyLO4mkHEeoNjBQPiQw2ZT3hgsw8yb
HVxpJl75ONlLZQoC5yyOWnDnvpS6MwbLXCp6xu3zp+Cw/VkkVKLgztvUC+l41fmvfzoUPVgZ+/cA
7bYgbCxnO4H52vHdHidlTKw25M9EErOlxqd6TxBVOK1JbDDz/Lt1ULwZGliHaVjV8hVG2831rDDG
Zc+jomvH8ro+Qd/5sLX7sgoPZdTnE6yXCGogVD6ufM41jKm6gcOs8AlUXmSDMGfhJeO0e8LGgmGf
oXEuUeJXtFMKTdBMn1Y82cpG1GG9n7XIlZnZQPVXUpETdwdXB+b4HPvZQu3KgxcVF+aq9FfLbAsN
U4ppwlTO2Kb8Oqd2MWcPuPz526U/Z+kustZaL/v8tjTH4XZrd9UCov4HuWFzo1rnnp0w81W6N6ui
HbLjYfiFQodtiLkrI7i1Wv/Yl7ce+uI/UjeuFGjwfARxVNj3cxF8bR+C6+6WdSzJGSOUxjEA22eJ
aZfZ6WLElBwXV9bISHRq8Er4YoL5JkMzPbELrTpLxrowlN6sT2a6ISRMsub7j8WRWayBqGtY0uUG
tuevCwl9QcLBwzjp+DRrd1Hxm2KghwMXJQ5N1D0NycGNaaJMoV4SwIH8cNwXp4u6OCgFijN5c2d7
/3mMTocp2+ndhPL9Ti4XL/YaTuJJEI5sJiVQM39ie8C6n16QNdvgOTXypisf/zQq0oONqXhoMxeQ
QSgGgAnhdBGxTDEsziDpXVkpriCT2394YoqIoEGbrhYuy+5NPhoHFbJXfLqXldSL5Yo9M2pz2kRH
oaIwjGzvazcr3jGkYvzWyQR/gwHD+TqyknU8ByaBd4c/HKBnlwzBEl8nJxZ+uTCGCdufby+2YY3o
XAwETZG120v9+GKwSm8dM9xu80GYDSQfU0drQGECYPOffy0DSXKqO+fq+y0Y8RHHMQKBLaAGdZuW
DPvTWEjQ1JQR4VCHjrbCu3JAeE+wmtNq4Qho5JBziT2PuVn0R61D1H+H/gKTFjVV58rCLtp0tHuU
Cz0waGo6VwC2avIetQ3MF6MOyUKBlndKIYBAurtnF2lxqV+mWo8PVXm6RnxdQIk68lu7OMQsNdEM
A9umfTifPESK014oSSEBWOwMAdr/4v79e51VzLbMwIQKmFJISCDWVa0ddU9hmuHNrQvEMHs5+qwn
lDmVpkax0DN3s2LMVck07vyo5hsIQXOBWZ/Cp/WT2UbAqSzFudMjHH2/tUvd/Tk+5hPT1rtSOfmX
rI5L+l4LKPhIkxmA2AUnEgGwofd8N5jv+uGQBw9IcYyuzg5WMX372/DDf2qEebvEgunx8qF2dOOD
jgKCPYPxEM0DpyPn0Rxi5e63cbM6PQ7+kkaxz49fPS4UzFMRw4A7VFLyYnu8bNHNtRBlApx0i5yb
Lko/nFnySFIx3jUj3oZwF9f6TB016vjRnqp1IMNqaidZq0QDnGDZd+cepe9S34sUKqN7qJvUGq3c
xnOIYtQlMe6RZOowu2gQ0aNcZ5r04LCyF4XJ1/ZnxXtyW/fkUthVrFG+hhMMj77VjfqDohopO7Jo
nojrVOIB1EDZlkAvSm50aQu3yi2UP6HQprKxqz2Gz5/KxeBLbtaYUXNzoxHPNitKRoJXvd7xNm25
V6U1wroNga3Z55yIHcegZKiu9Ap6ouhfkobIHMe+LocEjrV3McdxzM9rFXQgxXqHWDYVRgfQlwcw
2iD6KL8bClRdhH8pxqciRiibhwCMbNaAxeMCRUhyxRKt3mNoMKnC59OYwcpoXKYgsCOJNvrLKUIs
hllGDIFg2Difzf8oaOATfU1J59DA0GuPZf/hv6lp4/mzD+9tvORPOE/zGLFHSk6GXPmjAyIovLl8
+I9Xpk96NV5sSeFI/OYD6Tk5S4/mwQajH9TsypTn4aPTNAa07980Tdr6qkWtReu0XyIqefBW0aWF
NH+MD/a8/vNgcV0piz5mHZpJKdDZ0t68Nhwn/aMsq6IhD1uAwW8MfDORYc800uVGicaYMuzDCHf1
76cZN6r5GlodV4gegH8wybO2xUbpY7N5gZpdLcJYY93gK7tnvVgKiweoAiNrjPtT0CZxbSGKA4uS
8uq7rPNjNJnjHHSUnTci/6gBylcCFkR0MhQF4SRF1dfnbaZmuJoxMG75Th0QYk+9C+rfvxJhs8Ld
voFDKhiHjl/NSUPsiHU6pz2d06ee4/aZNM1ArdwyzkQKhbiHYs3DgEq2foZe/3wqIeBwMPvM2wok
HKu0IBwcKAz7vMEsqEcwBhiWCXINHgEQSpary4k5wC7chIce1oINVzJrwmlLv+BszgrkuF5dtx8v
hCfq6/kYSlPnibzaM9zrOXaNW/Sp7/VHMMvSr8kqmx3LhWHVy90C1XL0RLq3sXV5YDpS4TEyQh3u
rdfRWPpDYee8L8WIeFLkCeUNGZPpbrPnB08Ot7bBirNx3qqPxIeoPwD0lZGAZGzuTrzkVEXAXBTi
Fz1oMFEWWoLnVsEdDm2ug/XcbJNgJamvqaCIMaT+iXT9dnP63+ZJ0TZy41B+Ng9tbQ3a0xc0XbdU
eoOnRrQWF8DCQqFdFVEoPbE2SvJ6h/fHz4c5DI7B2C6ffaXujEZRPexuLYeCzurOPLFW2rTXKVsK
zVlBs9fHwV7gLX5YqMO0cMdR31KtDU+uIWWmvfxlyG5Xh9V712TRgRDFycUQ7sbC2zCr3rRvknGd
louXnzhAVa7S3waMpNglLK3MD7Gc6Nxbd/CX/MuOIoJAhryaMtRTXqjPxB95nKu4P9UeH1zGKDf3
fId2OwTcdn/HLeY3PzbZ/uqZaF9WqXI/NyxTcy5/Tf8atlX+0xrWcIaIpQ5+QtiJb9nXKT4e/Zj7
zuwRZdlJYmUtQywecowilEw4aeh1QMLeU5a6f9sj4RQvNFq1T/6x+Jf1idxMdnw8yxzzrbEhEKBk
sbItJAvyj80MB2WbWZrxUkDVx4jBR22SH/4NAninvq5BQsLbkhEI7q32jvwrxRkObDZNsJiwu05E
J53EGvx+WMufeIAUxow1kkRMi7Jp6gZRN7AQKkWrFNqBMn7Rd30mJpMNBsC2QV8k+JOUAkn2tfg6
frb+l+PN10YIR6kwPRfg+YOalnAdXhmwZr72e2Biysuu6TitApZvD224LWHxXVp6Xc1X1G1bL/2v
29k2IVQyCuoXX9spJAXsZelEvG1DzZwcuyCF1rtba1SiOhlm5Go1gg2bEUxyRoGK8uK+HhXzaH3/
ExUk69ousdN4l0vcVl1KkEylonPqTTlUtmv9Q+hHr039YqztE3UJBHjemvxDEg1EtZCuxXRo123o
wK3jU/arcJf25CVi9Wp04OvNboXvDb0iOgUpyMVkeR5BHOMwbaZjJVNWGtUo09TPy2WFSxAk2F5C
nxAARGqNUOcdvXtIym715EatRd2B32ivsSIChHAtii7Pt9itQAajuxA8l6YiJwE+uI+PaL6M6Yjo
BMXQcpi73OW2x5upRGNEYbCMPpfMOCwI+ETjPAdy1ruSDr/zHtuq+hd7nslifI0HPKKessk5h5gS
OZbHX5ZKaLg5QHvEoozKSb1V05w9Dqu3+ZfQjQh9tmcTggNVYy+vjFSC9aw0LWhBkiOeUzklRbgA
28JApuYAeyV4UXQmTsb6fgaNOxWr90voYDOdY/qjbNld2p+h7osG4PMyoYr9G5NU3MQMxYfaKE9v
yZJgZL2cm/k7BmPhGb8d6erMxxAKhnlgqx73sW2zAPQfZlwYH/T1tHvvBmk5DXudwLvEqpdIQu/8
uNF8zdKeB04Uygke9KAWfRCq7VN/KNQnVcRNAL1fO6OxrpWUZwJPhkDXl45GZz8gztUz9t0W43Cs
yLmf7Lf/ShDbBnHOyBQrmECvhZtbSHa+0Df+kb5po6+AAIIhMy6UHNuflr/Dkls8hbNoE3hBZYUc
sTt0TCJl8jrtyE0mIMbkG753y8r7EbzGSE+3fREyLjLPAQz5ybMAjdjX29bVRRgc19tZzqoA6ZEk
L0M7ZaEa0GHOmL4OOU9rMXrV1KLt/dC5PPgmdEml+XjSHFV662MOObSr/USqJsWGc9SpFwFIiAEn
9B9n70gC6NdLHOBYDT9jj8+Z9FoR34jxQW4kwhM3XZsct/8FSYyBvkMapgAMYbNO89RvTPJbR7+s
nQgKR9BqP0GKyTA8elpy6792ZY129ymbu0q9CnUNQ1v8RZMfZEDIDeRd/WTcw9kTZ7Z61cgp3h0I
3W+srk8fxofOsbaQaqNslvRtUOxBRzLobbEfPr3dQyo8zoXeqUi5ftDUENsDscoOZF1vaeUKtaLL
RxtSgQyzbAP95b+iMvgR4ts2NDrHR7i1kKjsksNqOr0nzPOl9yvNuDA49bERQ6RNpWBrg4FF1G6F
GzLhMTt2h88sLlJQoW3DfHpqOxzkUJS2f/A+tTudkQYQJsovU0Z4mM4xgJQJVWSChaJapG/vm6/K
Y7nimWhBjpVufY31xq1w3dBj8kGiGu79V6r/Fo3pxtUFyCRPdvKe04l5XZK0S2h/dAEcXEFMzFSx
MfMOWcYCguutmID7+a6KWtEjjiIwWuBig8XunYNTmJp0NkJMJor4+2p7OTNVI5btFG+PEavPBUjS
s7m2WAFVdVICrQ0Pw5+JTjqpto0RxbLCNwHRThOeFl6Rg4vkjVe7RHNPrkL3N8XDgjT5NjHv+tvT
hJD3bTUPJyW9IIRif97h/mQlje95MtzFzs6JAn4GpavEXHNZdRM/5F6dNDoN/QEWVLoQAqzOkmgY
MO01ela2bzR6vBoqeEt1Bvho/yXDyydyKMILouLToG00C1UaIMatxOHC7S2MQEXJlR4YFHJbtZ9K
boKST5JcNVsXb8tfPd6qmM6+YRkqu0fugMlncqQaHrV7h6+aBAJR4Xueznfko8IHDeS//BP7knj3
yTrMcli6thmnAKZlPZ/xxsSGeJSa0j6/1dkHhANB9qlkD6idflRQReqZOTRPKD096cyEmlQVUlLH
Qm1938g/WNF99GXjdnT+p22geAgLwm/5vEnLZ8drPEaqvdtPNWnivRClDFtp1MGz1GjX60EJD9B1
z2sfr/LmUonOHNnN9wM7m6cTQWWzxiA4K3twIt2AuQlwQ2u4OyzDeR4Uu6Of4in/MC4/DLlskJrR
4aXkZhZEszM49AuGxycaB3N1Nha796+P3yJLfNIRkQPRQ1+PEorvi7dwxbsnWeu7CVBKSfQAkiWm
ur5PjtnUe0rjWjZirhJKtFB8VuIbr41h/bqAhItCJVtSIa8NP3t9tJ1TWrR9ZN73arMCmUXwcGCq
Wueg77L40qyFRhcgxQAYz2++FNoLdIz0vguYMMFxWheL1/qBM3CoU22ioMOEIEdNt7tefFP4DPXN
SVULk+R0xZ4zgqgJiRlEqwdlH0KHKz95nBTEER2Lcay6+2P2uZ7uceXkJhJpckOc37mBB/d5z5uq
FNhewvNWDPX2Hv+6x6GOGO07OchrvHdVRNLofHMLe2Z6mqkHwDVhGcAHEcEB7HFclYj0VssGzfbW
aTzxKQfqfMvCM3brAk2tfPHTsCjci0ov7FALiy35YcWHRLTINSPqW/HMQn8EkaSmNX3SvKVGNASH
Ws1qvKouxZMcKUIl919dqoLMD680QGZ1pyXXpGe0+I8n8qWQrWjAgHrSfNUuQIDhu/+0oWPAoq7B
0rE9KW6XgrPHfDLMyjcYnF2a9YEmoTvE6M01EiRX8HObYwH0WyqKKtiMQqLXpnWtMoPEFSTqooYf
5oTdzCkijJQ1qPtoY82G7XPLg5ik6y/fC3ekkLI2ej151H1eeUWbhgEEDB0I9yv6N/aF/FMidsKj
k5uV8hhdRfqlbyzlPTVbakUoyD/XjM7GsbsyY3ro1yMb9gjc8SWE5tWLphU2WMENjGrKDhSfFgLM
esJcX/o3YyjVAi5Npxgie+Y0U4K7jc4BwbgxAnkJIagmZjZdFuMboC1JGE3eoCn+HUq/aYSbLp2j
i/piyGZV7swHq8BnbN8M6l1jtynDdX2X2iKx0KyWwhmPdCzL2CxoP3+5/X+hiQhuEc0/FtZNonhJ
y81x3zkqpejE2DIpzfPSaHFLB4VZ0wu24Swd3JUs0yh7F/8yQIR/xmEIlvGiH8lGkaC3evt87DgR
22bqdjaX8sSYTCrDaNs1J56QxUgJcpQ3n3hA3c1DsPgA/W5gDWZWuMlpVlZ/QBaiakOFYf+opMR6
yvPkofrx1+7NJmoWCv41qjZ0onz8ThzWaHrnHh8lqzs/L5lSBXa+wypIi74LkBmAfIDdBIJZXe5H
xNJABLkTIPuhVuOS12eK2BnMVhkdqutciHfNENDiZLcI+zmHJkaK4AqkwOAv/1BiBet6P9I917Bq
KIboVhYuSk820lJCW5cABrPrTS7A0YnHjoUogzsWWp8WFy7ZA+LAQuYD5iSC/xcy2xJ2i5p50tWm
6Bt4JpLGKWkQoKKLVy+psn9b6TKJvyE49jxxAVZZY+q7yEAngkU+KXKuil5qpmM18htmpxSx0DvB
cJ1ATkjQSUhFUdVxtTZxVMkhUxzcGtLCkG7t8CuFqUZuIgel07173wbBOCclrXgIy/NnkisL0pD+
OJ6xPv9jKnMee92GB6rqTxNee3R66hNWUg1pYROe3f2Z2M2zy799LAp7DfCTg2ZROgGWKb5oGHnA
3zEtcFt2sPg6kosinBFFzJd9VkdoEKq8f5WPXuanHWP/0JhVZvtdt3IydhIr81i8awJ1sNxkTc0S
SZkeEOTjpD3EaWUKZrG63FdPn7XSCdEKrr+xHB9Do+ZfwuVLKz7L6rGBjXZ50Po70p/UgSdskBbG
n48p6yH/p4y9DLCPVr7+Iuw4/UX7ccqrBBdDM4l9mT7r0bIZEvDhkx5JONAqRcFyzpu+F8YxNsBQ
ViSCw2nlrBRWR5/7+esf61Y4dtUfvvlhnxFerWi1RIw4bBFOXEVdRKW3doIAnwIb6l8SCTS44FB4
rBCP78m8p5R4qDnRjIRh0y27+E7dd2evGM/Tg+8yz2mz0nSv1TWt2Xo0SSsYcbUzeplD93GEf+4W
kMO7c2p8tN3dWZMk+NbmMXDmAiEqBsLI39IZs5hJH88fxzV4OlXtJ5R5g2Us5V3aHuNWz8Xa35Y9
S1Zxfn83QEaVlXMegkP0AGvIrQvBbi3WfKs2OCM5mCfyYX3zSfYidxCjafuUF+ULVYb+gXC10jrt
sXKZIHE5vk+I5/Z0zQ6jpkujUzRGoEUOHAXkxyi3FHhgLoUMQzt36Y6Ef4GgLbxZyWquo4tesN1i
/cDhQEWTquvs8VJOmTcm8IDSReUBSyZxLRlALLbaVvC8TUFS9EaU07g+VwWPlqpN+4qnN96PaX0o
ARPR5npSEdvLCbKYaTX2ZGf5k7PFP6InuZAtfiq8iC96AxyAbXXFxakkuTk9OhLU3eYNZSQnQ7Pa
70Z4dL6Xz2kp83QNawKc13L/fzDnXdUplIOFsJlQoz3uHVcDBHPK0vpJE9YSR7AYHlzZfPDyGcHb
y4Qpitohwf7U1odsGB5Ix+JOKHkb/8FpZFP7+9ZA/RmHINQLcMRXGHP0whI7JmTkT0uaPk1g5PgG
x/IVvFKvgsRJuy9+cRV7fT4+NLSLZLlreE9qg/aq1qiHuPMkobCE/eu86q2w87XlnI+gAuFkEQfh
QfuJK49Rqfkx1VIIWE/eVlf9JnFPOx/4s7kn07ySHb7UnNHSX16+Gl/2oaD9f4zXhTgfYJbEbjfk
12gqH4qcphePKDVfX7dYi2+CZRL1j1EIEWjEVwVlCwLlQgGaaLMvUTdU1g60PfKMnQj+QgvOWLge
JxHqufiNhOBxYJ5efTyrvj1PG1tBa44MJSHKe+G+jLqefSVrEI6PGsRT1y4nGQih+9AAYW2PBiKx
VrKAFqipr16f9fzxerPujjEm14UZe70wt+8IEMk26JsAPuNqkoVJoAZBOfgy/PXlyOkZsvTsBwIq
0LQMw7na2fhGa66Axp/R6c27a/YOu1bgmRnwIKBJbfCWKKwyvlPbmPA/LusY3NlUFSaKuYDMPnqW
FAzqys7zA1Dj4qVXOsAQmIHnUMyLsCGhoPCI8G0f7JX4x8CIMIDLXXB1M9KlS5WiXYJEpNMgSRJQ
EBfJ8uUO9d2F2dqouHAFUUlN/eriBnqqClxvmihJ0NFH2+M6PafjIN3Lt8g3/hvgwtaCL1BdktjN
SNN7CDNk7Q3xC6uezPGxfOUecNdVHZ9B8fQfcORA13BHmSKDdIDQX4QGjb3dvejozknhTaoMPp0o
g5gKsK3u3FvQH96Tb3wxdwHAMZF8r/SjTwvwF1CXk/w8o9sU+eAK2pKQreyvlPgdfb2cMPbERZU0
dq4vgbLGBrD4eeL5GHKsCsNznyXDXZZCmMirbwWjWYkEYcyDU1LHQ25EytNnmWjReXWV3Lt0JIWu
4DhEDnw200aiNeN6saXKR66BMOTRn64I+Wgh6pmGR1jo4GZQSleJnY5uKQY2hzu+/SSnqBBtwU/B
tRsmLmf399h1f/jGd+kulFeycXyGbPSK2u1dy9naq3yQoGrh3pOaf86Txz2FSR9h1MzduwOlg9Hf
w7kDt6EFKGFI7L+EcfHip63gFYp2poZaNB3Z+NlbEqT/ovG2760PLL2yIgktnokkT2mXzKoMOQyr
Wpy+EhOdQJwWDSSzuwu+zNhRi4Euw/F1HY0nbSL3Nb9E2zJ1VDIkhO0i/x0pA+mCx8kydZXD0Jtf
6KnqXcLxinWv8GWmJ4/Pllg1YjlwPa+XjpbBSWQbuLBli4OSO64V2Bfcg1lJdmVeKx2uAaYzKNX4
Qc4l9mZiX8RDkH4m15o548QA4dD6oaF8pUpslRRoyW5uPy+6HEEWcYln19/n/dO2lUagwKhW+2zw
DoiSKnx7EwfYHDhpxyDBzAZvaJ1hFiEXfgTQfQ+Em/DG2DvT81+8putuSbtYr4IyKdzYLjTnVHF7
CywJ3DAekibgb1PEZXlpLw+n2RpIhq/Db2KVIvoH/5O+AlbMT3Njcv+4r/zRI7BFrhB2EhqaJETh
uqS4XzLF0qo4lIw6+gM2+7wsKYb21R4/GhsveVvOddwFCtxEhjrkTvYtWJANN6JfKlAn0nfFA3DD
E8QigsqpHpkQHJk/QLoRFowCLSIe6r7KbdKJ9GBc83s+TGAnhOKFvnw7tKacg3Lkw+SS+/0kBqR3
HbDUgPsFgw4MM7qy+XAIRQ2Zm2rWfBeBB9ok9HsgAX7bKk848hvJxWrYCRgypa1iO535NI9HMvQr
Sc75LbxmrQGP6mJRF8aD2tw9KDYi07/ISV32q4yu6Vj/K7ewQC2ntfivyu1BzKA5Qa1y2VDsM9oD
x2f7KVJ3AdlUDUDbRUtRDmoQu4/6+WfdEjgCCRBdh7ABiErdfd6vDmio/o6yhN6IltQaQCfu9Ura
intJgBLIgteBreNr+IWYkEzU67ma4u3/x0a0az752eY+znt11CNOkiCbzCsRT03Kx+13e9LRIcXI
kZy/2glb7U8wVWQgNVlrQZa+W65CgHoBZ5XmUBXLqHpD4+f+3ewc+BAloAM9yMrxvDvPmk+AEKhg
3zlH4Milw0eVQ4R+Fd7dxWbmh3y1DNFrWPhNjrew4sTlus09NT+yIvFqt3XP2K1MN4SXmpp6g14P
CghEzvJrA6AsADNGRrgknrmxN4u85DEtA/4Yk2K54cylVr6FKa1JYYqKEiaUsIRA0m5KpH9YIT1/
OpjX61zjvopRk/P38BicrZ90+M9cCgDuPQ7mux/C+bYctTeH255jMEkk/KG93LumDAc+FmI/WbNk
NtyMA2rDfyGvCISpblwx5teaOgZOHx4zLroX9Rv0UqWGuSpmtB4Dq2cCZLT8LqWCeovH+bLeAvcF
VkXfVAyZ3qoiw82rrcVLMcPmpWl5NZ+H9JJwI3e5yP1/yG+/dODhjM0SUDaxj64yynxmZdir3hoi
r/IgJNvtjG5X6DCRhr1hNZV13qoMjlfq0Al7YaBxtolPS5QTRuicD1B01/eUcMm6t/ujhGuVe8Ua
VE4YB3Re+i08NSV0IaDZdTAhO8SilciXZLFmLFYt/LVD7hyIUOdHMFnY8WucRBrdFWby0IxGVmCb
7mzIcuq/bxOlp25tzxeJm9ZyR1zDbXGnbCOHBz7/N05AlSnj9JnizFsyvZStG0eTu1+9WTgUwsHc
ll2T9Ot2/CxNYPwQpP694Oi48H5SCwJzaO5JnPacxa1Q9cbYbDU64bxsZRPtFVvYFcOkcIkXGewD
f0OgN8eZ4fm7agat9/wGTy5r+m6J/7Rcvg3UqBavbV7IGbVXJwncJjHamPtiedujyDqyoYmlWNl/
b/QRNIWwcu3+KqGHanmDmxLtQCG9ekpQl73YYyTKnvsBwfw9Jr8inRqxT9n+sdTYK6d1uO3qrPEt
AMILLJ7T0MCUAi7/xa+jc2R3S25+wuoNawuPcfYekOymDzyrTy2JsQkxYP4JenhKpIcdSI6aH94D
tt/rbTUy4vgqDBScwP9hrVgP7K1vtP3PAfua1lvbHdW740q1ZfVr/vrqapIxIvQffmNhwUS3e8Kg
9uh3DcIHLDSfO4tkPZaE5quPiBMrK+ZYYPFAUKAMD/9Agh/c412DxeLKu/iG7qFPchTJ/7YVCO7w
SK9U7AktSV1QoftDz6zGhvbRFBZEZciYyStl7pZai8qzDzcCGE/P+rVMM87Kwld8bvOjR+GNEV/d
PghEOMbJV2yUzauLbicrKmdc3H2u7rrV0xvf5UD0oHex1CvlJooJn+SqRgyBq3YXv/0a+bfwkcjh
TDGlfbZ037RBpuGTvswzWOg7MW7MBxk/QpQPoHc4mPx5ZLyFySdSd6oDwce9BpRwSXbUjHIyNv7g
H2kKAFTSZ/zqKcFEyW9gGIE1GkhYLzan930bCm0+ZRrwq9JxVHcoXFrsnZ5a00G0JCWpspS/3stI
T/0d3+pgmBBqc/ZlbCKa2Xftb2PvfozXDAN7no6CGvo2MSqrzf/uWozeFPqyHccuO7Z5EvGvLqvf
El+6GaSvJcy4rP9xbNM+9oGAtRkTWbDGiy23Q5t5871g+4wMLIm6HwWckMdzIHOIjE62IUR65ipX
Zs8EwOAhSrgmOpmkxWYGRnDnz6scQaB8GpbYbO7mE0vRJ4HsuS0DZt4EP6vo1/wf2BliUooR9Bgy
jO0B/gRUJNj1wcvzWxju3YXpjPBc4bEqTD7M614FwoNqyzgt1LqwPviPdWSnAQNqDxBFHWUjD4nn
+yGBT6iiJcVR0+HlhRzXDkPlTbjLMdpEJ2IzdbQkxsn0p2I9X88DntlyMN4MoQiWKbqa4vN7C/nr
AT+zqB6h+rKqpbGMaZFR+WCyj3yBvro0bBIEvLib5d2nbMcnnvZujT4fqL/QLmBcqj5ehSnxwiuY
+lvCHQ12gNNKBPKoVkQuZ8vr2LogpC0Gn/TO06MP+LhBqigHq5v9b9zkm9/KwVREL9W0mJdrj4Qy
AMOCo6cZN0khhEr+wY6eq9jRPd8THxdRQzNgUj2InYx8/lhLkCjUzlBNVNiC1t3+JF/gXehAgXHa
n3MhK8rxGs1eHOQ3h6G8y2Jdmlbe5CfZTsbPZIaEUv7NJ0lZV1S/EzkD6ZkOdJvgijfXrapEwK1Y
Z5IFGQIqW0o9b12opaTODuIrfS4WdDcPZxBEyKKAaBOW298Hg2YIcJoRK8jtL3ERK9KuL740lijy
DkUR4gSsa5PzaH54b87vDT470iAMpWoYwFLCJItKNP2boj/q4fqup2xpNnEuPErxGJrhG0M8dwLa
xjPnlD+W/EWA+6d8L+Esq3OrZwGyWPf+hCUDr03UTbhU/+6JKYAZ1H2tqclk8yULKpGCG0mY8yE3
8xNVDfvSfDop1OYp6+jr0nEYIZ8w5Dh0TQ9jZL4kOK8y9WRFDjsqToa8NHcIWACjNlPDnIzhmU9o
d2gWrAGLgvjEOEaoHtMns1fy7KzQLRSjGV6xgYePQMKolaIMgbfXsMkepqJF2LScfA8I9ZjwJewc
QclH+ISinDmBIoDM+lHhfoGnrrruTaMHIW06dFlkCiOSKbqiYenSaPiGuzoGhm1S0qKcsoZ1hGlI
XAqDRSXmHPjc0AIo3KeYcG/Q7MAUfT3KgzN91FlmCvzwgMBruiGeINBGSCPPM/9JFmvXTE+rq9hT
Ha90FNTKpOThDnEB6JKdja9oC3+p1ICBWcc5mrYZ1+VeZbz6wpaoh43ugYZ23DWePAADWk83nSSf
DSmc0YWGQ6ejXFBXm9vc7HpCKDSqc55RL+l0QLxpT3IOaAvlOOXqopLO8CSKYOAPciBMndp8fRZm
lpgI7KDC/mBV1FIOQo8RSLUVjGaGCTzrYmWARSLRxtdYjnBkiOCVVFwakoH6fj36qdCwbgJf0lAo
VBO7xI5hdWp+EbXXGMr1fBIxQnjY7WA55+Y1OyfI67pjdz4sAoLrCVDePhJbOTA1MUKg546Z/6pZ
6Agdyz2pzjNjvLgxfOIxuNWa+uTJwtD6QIOC1R2ZWxY/JUmyCUpJQE80+gzu4eYGwjgHC5MY8H27
+ibWgPsoAnebfCN7IwO7A93Y1CUqCK/CsPLXfEP9KK12nuGCpTpTd81Bo8stHTd5Dl0iB3NCIURN
mO62jVMQExr86nD6/HcFj9/05tNQ+CWM3eopFTvEBvQXhE8TroYOVE3f2kZgr+HmQFtpgtdxFPUW
O49lBwc5RDHadklxFvCoA+IkzBKtDSX9lXzPAt+2B1VUlutrUzMF5c2Hh+W02z6a1XgNPnOLKpjV
OyTpH9f5F7LtMFnP//P1iVRLtjim/LK+2vOvQc2JG7JdRkhcFvH+s4FRYEa0g6W3IjxR44NFMFYp
RIJoKui5HQPu9lKu47oVH3LrP7upj6vnyan1w11VhdCHiLsC42RXwbyG4+XKKP04mycgUoUU0IcQ
/kGdvarz9PW5AKu37+BJB6JEVpgD3kZmSNexDNbrHfeRAwPeT87HrMcMNaQ8rSMHwx86Kq4z0PzF
8W9eSUTaYediC1aJtQW/XdayXlzp0HExzXgFBO1WPBSLzwJ0yyJvNVI2/ySy2ushh6s1BqshUtIh
SRbwTUqmo0zzHfQzK4NbQZuOfQDzA2krMPOlqbnXPr/ncXktrkl5h1N6JejRskG03PVHPg9xJ12p
MGZv9OPshGn1j2mrgSlPyTyNnAmRKSVGtuJQdn+niDED5S2uHWCJ4e0NRS5MIMiVuXqCTZ2PUGW6
TYP3avTIMd3WYERVNTFURuIpuL51tc6/PhEKs41tVemezYVVVG/vuFZw0yaj86XKG8VKX3W8kH0d
WJbC9G/nezDyLCIT0qo/ikCFKDEZfhA2nVpZwIRkI9I+IM3DROBIMrqCfDsfG51Jny/FZNaReuyX
d4u+xpw63yfmqSWNz6mh2TyogL4m+1erlux6z4oxo1Usg5Pu7Q8+yBQ2RAXaTNF56mBP65blcx4o
03V6qqyzLmadn2klo+ko5v/VHY84tLlrf7iHRdG91DsBSQSgkJt2AdpMtlyUPJvMh+MgIXtqxw/n
pXhbZlYIkztGwlzr7fcg+LI/XxtQiehVFaTsnLAHssLViT1Vmoq8KYs6zVuMA30kir/DeEw69FCu
CX61mUtPHjAGpZ7Wx1cunjJpmDfS79qFXk538TF8IZkCkth0FTokWIrvmk1Egd6iTBxVA2NZMQfs
9HIPjUA2T1LBHLi6sgzKtKSFdBL/H1qGgmXVf23w9SMJ1CDaqVNsB7JqT3tHtNx/wN0PAqYWFwtN
br/FSldnoSwx8dkZOw2R3LU11EfYhRW1p6fQwmiOTK8wg9x6Tzof/TwLE5YswS/dScgHJ6Q0Jwci
OEnuacr6s706ZQ69wIIw5sc2cLJCRFSAkEItr1IoLEeMDzavZsnS3h8QdR1x83ZdEvkV5qxPmewq
Ty0hsFzH4ENLEwep5MpC0Wvx6PLeh/2Ilaie5QinqN2qppCxPJW0sN5MLZ0602vJCyRwcbWi1q1e
2z1NYrDOHdzq7Su5q4S7s9RrvFuCv8dI2FLvOMQx/PAk+F931DFJCryo78rAJrPWLpDc1P3Ztol7
CGjUxrqSc63att5CRB7JbLP8hGfO9UQrCzPEm08ef5HoYB6yIcujJJ1POm77xPOzjHZ3h+Uh5b1G
X9DGOSZa574+UlkyXMkd39e87D8wWAOFB7WIkJJ68vCcR+Rym+ZEqMJ1WeynYm6AXCX8PkNp0Src
JntNbxlR9vcR34LUo5aiOOMhxHBHU+bq6OuP5CXTqcVVPprLXyZY5uXRAYbpSMe+cMt8E6Oze/F0
eF66JePE6jGvrBzmnbErWBasOZg8vghcthRMH5XSu4w8zzwJtYX28h0t6dxmSuBiINRjzyZ6ciXX
lFn2XB7JBRem3f44tvWV2SyNRuBv45vkvLFvQ2Us4UbjuOw9odwwcVyPoi/t17v5wN6QwiHzJCY9
O9tczS59M38bCDVXwMVvHiZZWFEvF2RT8qPrS0SyGoj1cACA6sgDeiEOdGB5Li6IXiUtL+eJ/+Hj
XW87E3ePviQC/wpT0b2LVJTvNxjYAPOXWw2jLhW5tlUzOexL+CrFlKH2d0jgaBtcvRlt+8uAHZC4
4y+dwBx3RtbnSsr6NCY9OseU4rdcvLyg3Dujzf83gXsiGEgZqYpkaSA3dGZuTolZIXuoZfi/VEek
uf4iuI3cutyb3sgEwA5/tQX0bvIm4oBYNB0WIRM47ApHWyUzzefPdN8Exs0P5uvu4kW20Z2Eh+8N
lyUmC9vD7jERWln++DyKdbjF/gmfPfWChe9BPX8SqNOCuLg/UpEUciUgB0QWpf2PZX4G911ew4co
2afDTzaPwV+tHqUgJWxzsxsPAAmjlFMcL4VCPyxR8qR21RiS0mVhePaiyPV5kQnWz3mZcaE1p4IL
zdAMJIGWfDHLwnNQiCYf8dNjHjKLc4eKWWgPr7NEMt5lMwhlzw404e3cUWnjtqCX6+iC7Bwhgxx3
u5UzyrCkuifpA/71zU7MPP48VU8XK29vHxSgIw1V6GoOkHM3pzd9bfrSv3Wq+cYsBAWp7IoHDGRe
A0Y3B7WbQ3PmrZcnPepk9Ot92WShguHsEC8fDtzDfB0udO9aR9JMInQOGaXNrq4pAhfoEBKe3M26
/lYyNIhrPu7KxdRG2RJox4VRdEMNfB2lpaUDlhceU1Xcz/RVA602lp/VEg+dOQ8qrHCG0zUClTbR
XGr+yKi6H46ri4IkTDtRGTyFvJGWxAQ0WcVSIdR700ShRr6Mv4tQby6pGlJNA0NP7Wi/FRPMOG2L
+oyNZNcYRZN66TaHpZqTU3sfG/NDq2QQErP05+AnaKVzpbe/VTsef1CJIsnaKuAdxEmUUX4AcQW/
MPUlcWTW42UVuuz77ZfI0ouENe5GnL1sxCL4jELdo+8M7YyT16RWwibNuYmI3+exmnfiE+1E+W5l
6Acuf58pwSnzHMGxhT8XsG6+UDW8Bv1QvDaR0p07XhWguLP7kKuZQRbjiYg8q63FxCXZdNW34AHz
FbFAKXN6+Qjs46YJrivD+fn0tT1kk/zNvgNbEw9XNaYRwcZyprZi7RrBaam9URNU5aduZw5hgqbj
ZuZT9Lis2+jODI6WYTrOQRTMNXhSUpgkAcNn6iByQv4IK+IbaiBI7esA3wcBkLRN1XaCPm952nsP
b6VJt3+DOUmbNvgw2Bygo1FyIu57VB2+UboXIfN2Jnp9jOb+IxlyytDy6ED156TX+qBU5I0zBiuL
B+qhx+e/r7M5OII8GFYbc1fhUX7Ct+HuoySAZylB+ocS2iFTCd04hh5JMfZtVdTsZxqwXFDjcXpn
1XBRHn33sKSrBm3MAfkT7A2CmOfqJre/NJfcS3yBNhgd7NJ7WYQite+zPVbnEt1R62o6xSKFlzjX
m0DKcFG81b0Ag8HtmfG9LMEqSFUj60B3EIaf5MSed8ezs9abOzPlNdmMmjvx9Yn0Io2m9hqqjsh7
7EYAfCdPnZOHsm2tJGgp4iwAEl9Csdhl3Fl5FANUq4uFo4iHwhe8ZXDAchdREcAm4wngVtYodFYs
FQL38QXLYUV/cY3ODVwQW0O/NJctkCVc3eC9wcBYbXaWM1iVhdrc8l0nkF3YeQvXik4AmJIROyJH
IFEFWG9zQcxzNDW1VNTUL4hGhBxWnTIu8jsrNO+bOkvti2wzeq6Sdl1YQsuOZwO8VPcaInUwVmAF
r548aaFEtLlq9eV3pw7+Z83RIzD5bfTGUQc81lHF2mk1LH9JLcZmiplbuhLNA9aEbUkX7asKdYGm
mVOIsK4ukL4oJcdbQn7XoWKtE9C7SQkW9b6U30uvgmxAqO6i4kll1epbR+Fc6zXPho7Hfoaf64qY
6MvUxS1yhPXtz0abAIAuIc97xPzNvKCU/V5y4hbyZvSAmGBTthzBB+4O3YCv843BKN1Xh5OLxll1
fcryd0BnNhoSvXhd+OiwnTES9miv6v4Ig6Vj1QdfO+LMvs1vg19PhZenpoMT7Ah0ACqgAQWqIIAz
J+3StfyIAHn+LyS1Koa6TYS6lUknx3NlDxjvERvDbjW84uGzeTq7Evz+t44LxFPDzFGZHAzX2WLl
7FNlQDrtaMMuo4rF+c7WMVLfCEoFl328cbFhXjyDkF5MwbIUc98SynZdIOqEvQ/1JZ6E6UtblQjf
B8iufSZgQ68yHfIPj3w+A/JhNDH+mzQpuTFfO6SHRlKc+K6V90w+R6RF3ihfLX11vpvBUJqiDZ09
P08OtZgusFFbRpvFlo5Hzh9yDHk7tlhEJ/jV9VzRYXHWG9wk1xElTQGtK2LVf/QmImEVrlVJbMp8
chFMNzc5BdYNQ9YS7DroI7HPzlRPj7CJ5Gkhcm8NyPPK7rQ9w0d5YaDz9mRMcajzwuvSAWMfnUSZ
LNgXPKGIH+/46blOWYggo4N+3zRYxsPNM3ch2uZqMLPQPLby9gbk7VODBWQH3AIr3SbnajUdelh5
x12x+7AzXy/Ni961PN1iVvHyOr1m/FCigK9iNaT7Y0ejwHOOroF7mfkxjfRuC8sHkIw3ED8Bl2SS
t4sj5aKsbOVRvEuMQjykTRSOaZ6I60dHD3OPAQYLzfp3TyuALEX75qkERL0Yx076zyRwo3MgBgV6
o3dS7ShfvvS/PDk+xJYmmwzp+ltUTrDVEWqVvCrOQFawXzzWgZE0HspFl3Yp1w8IpTouA82k11AH
1aFosLtNgZedNPM78eXBiMVwsq1aGsCUlIfijRTFo+hZIzG58UwDG+ScToC7ATabTdkehJWw83DF
iKPRNwWqNcuPJm+m9WRYIwqvhqIA/2FI94krL1MmI3+xj2YCLh4w5UUB0i0O15F5riVBSpu6o7k4
bflVqKKLB7/XW/RxjK+nSwLDRqD0vQN5rTNU7lgk6O8IRx/We1zfUXnoCOJaWS1QCE59hBDBTmYn
lS26zEwoVWzyvquBbKpF1Io+RXSxM914a1cJFdHjaK7z8KYpUEb5jkfcet12TevN1+8FwgUk0k+f
FCPZdAAvrrPkDeFfQc5v2BgExTx9/IRpkRQqIUlB5scp11X8YTIv2APcJahUj1eRuuWDFYu32aRf
ebT4Uy/dIreEuT+PTXF/ZFIL19KAkzlRVDajo5Nx6DbqFKB/N8Mbp4ITVUloxQqa5tJbwrX631Tw
TlM2Opi8ncqSAuV49AFJeDK8INm64aKmjx3naVe8oxjiL/n6olR3Ft2o8ZNaIXAm44pvjNPvRhAV
Vyr8+f8xfQxkxfbKA7dy1et/Aspo/5lNMJzWliskGh7KzEynFohC5HZcmWx7Cc+gVym7n/R60j2b
X0uau5uS2PTID2p+kuQcElP5he5lSUS6VCZb9R1H4CjMUrnHm1zlvfMSHb4VOtsJRDeUDgl7T1oQ
8/MzskWHhw86fp+Se5E8TVlZ2ZlZIgwwsPNUQJWHhySgz4AJ+MnodPhZpE5GrIxdfH/TvcNqyNAP
gAXnk+eJ2gtLQqKi6VdwiJRszj8isUEk7VfsmD8MhU0XN3N2Ao5AUQcw9IpEZSsLCrFau+xCKlby
MODMdPBmBOhP1aG1bZq2JNNCSKNrj2Ju2olpcRtNIiaYhf12wJ2vVPX3NH++OA767Tz9ZLA30m7l
T+c3Gan/k3F6hbLjSVjTUd2t0vJv+9EXYXWzk3WiDyEKcBAM2hqR/kG89lsCiHExfY0+y6KIFql5
dvFivz7zzeA22B3zL84hHeJJXEZPN7PeNc0f6MLp2VARDAaaJlRe/hM7s+gv6p2hwBtUvNeYYnRF
qoGn1nPAd+zKkjFDoygCcl/y8uJkyc9+p5AqG7zKY3X06/PIKOtn/zO7+Jm8YKHYuE5fPlcOkvpo
fE7so8/aoDkDReBcNw4hLRoRqruW+xsNNsFhd+enCKK7GlVoAJki4RdmtD5jxpK3cw/PDPUAJ3GW
/fPP8SEaJ0Yy4+43u8o47Xwz046ymFae5nLqG1YkQQs2aeG3LC4SKcfUIuXjabjnEDTrfUc9a9Fo
0+31jXEhKsZKSs/101tvHcE30JR9LEXX/yX0kS68Q1rmUkWFO+SjrSFQ0PpZBMYCXFBg/XUBUSN6
QahxiE6x/O2M4TQ49T5xW5m0rV8GaRhZshtEz9gYZAz1q69mXCenOitGYILHTi5x6dUsvBA5Q5xR
fD3RAXKkJhOqYeoKH378Kl+ffSpXe3qyFcewLhfD7D42835OimKBgzuLcjk06kge3+JXLimyRpzJ
09uD7J8nIUdccNcADTDh8524EsiLRS1aNbA4YlnXGm0PGQfWdz7Sco7D2HlvAcnIvpVhwo9e1z7U
jSaX8YMPiAdf6EPM+4xyAt1pZ5vZ7p6vCTzCZPj2/O4fI2FwM8WV7lWO5AdKKtKVtRLBAas4Fzql
MPJdk7UgyYRHY439pWIonZemb9qwrwONa1X0w+OrvvrDKaFJNQUiUMVZlBsml2IdykXHbOJPDbfj
otdRKOJamdIEwjzESeA1C7LpfuriTkVLZ2QR5VFPDPY5sqCpOL5mUOkGdsushoVwh2n8PHH2oE+e
h+BWj3MXj3jKPN+RV6dEfHHskUwxaESetr640cYvQg4kfPkB9yzFXRL8WmS3bpwwd7EaLXyIysyv
V9rU5U5cdWEvzs0nj9Sz3ddulCqvw5DHcGnLQZgfql09rCpKF0CT5Q1j6W8vHcwrMonarb4Wy5Lq
2QkBfC+QXm33/NWZ2LuwpEnUfXyvUabokmrRq5UTLRNz5dQgUSEJpA+jmMagx4ctbuJqpcMsoVMU
APMQSv6uiaR7ZrcjmiXn0i67FIJrmuQILgjlC0w2Pv0Ut8lQh30o+XLUAqyev/8bUhQfRcuhrcJJ
jCCSUyf7aPAm/RQJyqbyJDuf3KZLGwXrtpgRlKb/HsqioScO3fGch2NvjmQSgBf622rt8N4pPHnf
V1EuGdTpqI240XEFUme8BHJSypgbUy1SFbwH2ge4isuFFrxHfXl12k7ni/8sFSTG2KTohCLHvvJn
XdByx/1bFmCYJk1YNr9mqVlMFBhgs0SilZbCrhe4dRMfhWVMDWnPR5rQTLqXtPrRdicQmR+6U7sc
lciDnsxhbQk511szEn/sNmfR9i/rmXnPN1kndnNMmmj8g3WkFvjSQexBUEio9apmtjAFQUSGc4QB
ZTju9YoNReFfWS5N8HCePUOhtj4VN3Ewn0RigjzAjCZYgFC2EKjYuKmQjT9OvS1WCY+rga3SrOSo
W64ljtzyffv3nlWwkCk/34Cmh8QOctzTi0UyZuaxuJCKBOxne4KNQ0kwWZUneV+siMVoBRbr8Qfr
7ARAXTb2Myx9TgY7P1jISPgIJiol2fGjcTsVCScOIKrzR58RrKwEA7e0G5Lo5Zn1Iq2Wrc8izJJp
UYPwHejFQo6jkgPDswaakSSYSSb4XAQnRZ/C42WJvXXWjBvXJquQ2cr9Y6OrzaQ81zjIrn/iei/I
b2bstPrSneXjua+apC/0JgmQ9w0bfHmekHbn4LGSAA8JzqQ1tZ63nVV6JZ8PC8i+BuRi4vxNCVJf
Ax3/168DMrzehEj/1O0ZzrRcyDcMStTE+HJxaHZ8Ajfwp2E6eSSfvn4saDWxlkcG7fi2hFC8lBmp
mb3d5q5f44hnSGElhjxpdpl101iYcQRMuEGcoesmNCrtpMlkyIPXukIHT5pzsA05/4MGMD4X1jHC
+KWHKr1sIjwFUtU/0O3gk+klaPE8zFL+t5P+tnl2/HsfNx9A7lrd1Ai8paXPo3j91A4gQDVz6Ql+
m8p96NHnH9iFm6k4LSHvtRcpt8WKiRybryl3w7O/9xvHxriYz98h11MNgicV2zRJBxygtBAMwrzv
jacIGoy5CV7cYsmYEd1JiJQU/LCVmhlXYdbbXjJRDV+/Koh58JI6x6pb0bbVyvuzF8r0Go8Nvugw
zUTC6a7JRJovKSBUNXRBq9SsDSo+OzNLLJthYg01RsYTravvJ6O0of/6WEySJ9qnp7bKCwe8JKB0
GYBLjC8ffAaK0lRvrDFRCwh3Md+6HgAKf4y95xI8YKuNoawOjQIn5J6OGmSwRgWhMWAwJMxS69a5
ziw0N/CSqByN+ONxF6nEs/tk0/JPNbbKNtnQ6XOImIKVEBl7nyg4L3tHlJkE0AK+guBsBIL5FJDZ
YyuS9FehjjYrQM139iIx01YNKQb6UMKr3e289vNSOQSxO1uu79kCncVjWkfC5sat83vJW2kIhwzf
I83HnSlTeAUXMoJEUbFZ6QSGwd8zc2ktaqhj/qzZWvcQcnJ0YtKGKo4TjXcx5Cou/GUc9VeJKAbm
k1yFyf316zIMhhjf1+Lr4u53Evimjl9wdzAoF0ZQ0sxTcLMO1L5++RFraX4rZpspqOjYgg0z/nrP
ZcKRk41Taht9Xp9NaHTT0X5uEGJBGrjOkJPnThEZfE5CcZ6uUI84qsireZc3nS/58miL4Q1mCRwB
dtdwbbJFF7EojeqJmQLhewMiccrRxVsc4v2NUq1pmr///nYmQAmewX/bx4VboHouGr7vu7Uw8gWB
2L5VAl/Cv2KCJjYHLa19tQmwYdu8LbX1fLVaAwb4+imitKYSuEZ/LujjnK7+xe0EVtBB1sUE08SX
RsIiVB314eyM1Uy0Hr+N0ugWDl/wuKvqyXXZDKxRms1Mvh79gIO2biM2cLj9eQ5RCbIgaYPoO4zB
S0mJ5N/ns4tMaz1wUzMZ2sJzoWYvo4jMpP0OuaAT3P/0mMzCVSZh8mNykq1j+/FzCaMWt0wZCYWN
93tDxrK9CfT7ccBkE5VxX+h7fjJ23v/4U/+k7PfxVJjucHm2s56Bqv8qeaztMSqt0EqOO0hxkHtL
rsd9+VogBfl6ONMZ01c3jScpCHOQW2f3yy8sIALsTnZh4uFqFpxls4zlexED7kljnZUDcefxh8Jz
1+g4hafDUG5TTAz4NK/Kpw1JJAFewpo3j4phmC3MWEhipDhe7k7sd9xxW9abb6wpEF26UxS7QX2/
poZNT/mOGvbpydKaT3MFuqyTwEa8nynsGkHWxGp2lRGtZ+vy1n/lkLqgV8xBiVzw5tHSr6mGduZP
SYmEmKgW8MCv79tFUqmwBFw9wIhjyLEBG6DEJPzGkxov2jSvbWOAzzAU/HWf2rVO9GYWVbeTnFJq
Sm5uhnaz+M7IlzHdDyNFJb4B6elIbM+IudPfwxwkTLRwvfoopg8EKFtKsh0DhHSUTi4sYqhJqy+q
NgfuqpNR7O8dx8mbBgSeMl4zwuVpOKBVJesdXd+7My9BE9dRr7r1CffhZjYGJ2hVIkl21H+wOJWa
8aYRYcU4Ce+ZG9Mu0xFO/usI4U1tZd1KU8Kttb5NXB/BFf94l8hRJwfqIiPYwi322H6VZH0Q+SOG
i/cK8+RZ02WcFIF6RrcCq5bcHsul745AvrkdcZ0+o0wTrqqACk5gvX9frYB2Y6+iXubM+4o7Vist
GomWut/KXJm0b6unC8uVeXlOasni/XPPQoXMMGXqvuYgyUMSHvtChOoFp1X8VC7OPD+ijhMIWpln
cPh3WzM+Ejiy4BONydcepGD6Ch5IHgsSmuSEXaEB6BFMfKDpI9WyeTf5M1WiddepdW32q//UzhiB
+zSgteZWuRm7IdrxV9dyxaZWPjPXpHI/O1eZQidNZeCI6flv2J7o/gqKUj1Duea2iEV8elZ58+JY
pUa+6P4IMBm+dZtI1EPDOpFvtCKFyCQZa8rWPZvmisJriMwIeQZON84fl/QEPnn9m7hIZc+h6U2f
GYLFp2Z5rr7tUVx6lA0oXoTAvEfDiVm025+zqnf4pK1ip7YeX2EtYklrhlOx60zMc6pfQg2U32lC
10J70q1i1xnN+TrTLnU7Alr00mrzWtB/llX9b6kaNXC3VSxgQL5pQ+eZKc/IwhjkfPiXHd4VMWMC
JBeyN0FoW7x5aM9VN6McGU4aVvFNLFi0QTgWPiNgzHyNMGYAwu3NC3d9XPLXgVnc8/iPs0erx6zv
wyBkMpgWZwpLCU7ttSwf+uAl8Z/NkYnZ08D6IGJb+kmJQSpS8jCajutt2VLFCS7f/ZAGKb90eC0/
PlmbIbifOI2esg5IqJl8eZ8r5Wm2gNDgN5r2BBCN1Sy4wwXdkqOt57gwAttNgui3WawyO4OXcXuE
0Kh5epyJYrROOoWn7lwX28X5/koh/QJIub+Hwp4QA83v1tTMoq83weV/Rd5X0zhZHcLn2qwTp4p5
y4mbruZjd7uF6RRqOtGIPculSlUSfw2iuGjMY5Y5iIM8bwwacERCrTOg+CupOavzLwoTQnV5S9DM
6NWKLUm6TIQQfw8lmS14ELDVLNewfsf3ck6wRRZK+eJeIWVJDvIsZ6pXLVVioBHEJEpnbx9vqhyo
LxOM3qqvYyKDr5I/sLZGwZA4e/vJaDnmYPJfWxV9hwUJDgSj6DrmzCmfw0h6dpQZ4nRgRzNOQu4a
FmUwTIl8KFU0Yik2tbyTaUtlsBDqIOrb2WiKMgAIEYX+e3x2W5azOIqkKp4UqZ0U4+aKb//yu2I3
pyoZ+DGXQROzJNARCPoeBVp63zbJVmuqIZ3IPO0aGDxT28XknkZJ8+Kj/CR5YR2Tm8/QkQFqIqz9
kKdZxuH/IoFpzeNqfNuETI8/MU5ebDtbyHxAib3CceZfp80hK5ZsHeVOcywVNVL9JGx2f63j12y/
fFl8t/5S/w62jJrH52zY68Bq6W8ZwAr5S7tF6yJl8NoDN568Pc4zo1HHmy0CC2u2CALWNfTAmXxO
2pkI0vBalb7p+lyG6vxb+YNn6ek3UjoYABO6Stxt6HCz66xQ6qL3m6JLtzIDyyfC0J7WFlGrjZaW
0eC//u4mVqw9olFzFLJOEQp4E+sZAXcSEsZpQ+M0BzdSH8UhzPqVpLKdmn3sJNPVEdz7/PDl9Ozg
t3fv8G+PCQ/RZvRJIJRxrDBuh5icV2bs9f5Q0jNDxee5zYWsesgbXULWgvq5uUhvYfUj5K+0gyKW
gXRAip+VEzW1/TmBVuIjPEBCxT4gVURtD22zgOvil+ARUmmi4DNyIXdWdmnRMy7oddmk46wvGAQ/
vMx/qGmfDV/XX1/x12f/enx0AqQGLMERJekLwtClGBsgAOpI3O1neeWbRCAXz36czyexc8pBtJxy
t3dGuhedOrkucm3OPhVuh5ioQtwW07vEL6rcQGSa3gJKoyyiid12VcvhJen7WYHj5R9JRXugzLpN
dPz40cmOMFw6Kz8XCccsa/UD41Z3QjUVbc7RYP5ixqvClJG9B9qj8CFPTTKeO76cMaDJZ5yLzf6a
finAwL4pxJfcNRsl+Fv8ealj+jv68NkLDYKycUN9d6fn8clTIlbkXzXVRUY6//axrParwsZ9B0L0
GN0pOn7pm3ayRFlEvZdZmabFu1COVnkTwyh8aSg6dLpgp9IuyyPCZ6KRIlj1nbg1T+GhMTFf2oPH
IqSAvn8EMoQ6XULKdrQ31wEnPtAbX4yljlMyZU9XEr//CdC6XbbIjPTcu+i8av6eeUSVPPzw83Ah
HYp+2S/sauPmuAwRoytmTBFnavFcozS8sBODJfFZ7/uaUgJ3hLCtYw5oOleRJC9ivok9EHKFRBSx
eC1EgNA785RGQyE3OT7vt4AMVIfku4xBBSYfjMd3vHQSCL2ohQX3YPBvK9iakT1iSj22SjxBHnAX
S4NtVC4kBfswwpvUI+3vBwUezz9kIVy9ptsyz899/mdCLhCvl/ravj5CfW8ykRW9UlxK6AZ4Agz9
UqVsoeclqjn6dzMgHtZ5xxtq12wg9GcWxVpLLQXhFzIag7kU66EYs230T0LuPMwvvXUpquL/19v4
kYQB9BZ/cBmnDwnEref00+ImW3tFwQ35Wbyq/Y2iHB9PmJGX2HaXLL/+V+ZCdp2OTgGzlLzx5O66
gxdnutvu5xxSjL08jT1Gyj9iWsEQIG1uGStn1fhzyqi5fCaM83Svq+O7JbyIwQajDP9u0ESI3Mbt
eWJyyvJXiTCdLAIvPrKblErex1NvTXgWJNjxh00ecWiP3wYxMTn/m10+Rw8sob+E0GTBPgMgdDHU
1+xxsKmPFhlujo/umEWroxZ+h/h4EeML5/uXyf6wqAUiYItANESTFHbkNgpVEydEmtnjd9Q7PlFd
u21uJRvRwDaTpIdFbSKNln9Mka2j7W+p59qq+vSS5813RXAta9oPbFGaFqwIFoJtmzy7owxX062B
dq8ovpbKtyt23oFqPjfDqwCwhzRdNwuU5CIT7nyI+AqA7puQo3SAYjH2uEsOxYkqKDcBLElE0nTL
IbkSs02VxgHD8OXZRm7rgzqgL6Wa0U3S9Zfi5GGEOsGNajRLank1adMFRsIMxtyYqBYy+DGggNAW
qgy+egmx7fH441fn95MmPwwPf6fgyxgxCl8rYBISGGtYjpCUBzRep9ly7s9mnqPiEesGL/IExdvU
txtpzOPNO3ZkyfKkUlFZzkzRgSvuURyOnZ64+punTY3ZCtXLoBtIpC+Qo0kRxn7W0ACRkFXZkoqa
M1RECP/4YouSoYtq54F5CkSnV6vWpeHxviwI4N/MHIRf8fLme1oTLk5gNxxJv4bvl4ZHuc9vCU77
Qi1FbmVU6qZIs0jA+dh9lbBsasOhNm2tkJzQhpx28SiOQuLEK+K6iSzLH351fhDDTK7llKorSvEw
JCuqj5qDvR6h6cu4nAtu5awVA7jmznVrEatTzdiSjYqQjCLVsYgpytLOp8+/Zq3+Xk4BOFnUhPsi
fPi+uNquy7bmNSxLRI4Mhf0Y/veofri8SaCZEXd2+JwZAuHQkhSdSrdtQbFq5IW1yp/DrNkB/Hgq
O7STR8yEvmYomVWkR7GJuz8SSNbH7uyZfcQMXBqrISB62vBg/X79ZCenrMvjUjUCnAp4uHN3Q0jP
HiSH3iyHm8fNcdJtir76p02QhqkfAMpIfvoE4KWwwaPFTHDdPf2ob0WMpuUsCbsBK6D3BJV5Kkee
3tp2sVNp1gnhVwWL3NWEZbVWQYPh2Hp9fcY5ZcC/jXgaK4BpGutAaGaDg4PLjbKcy7CqhxQW9ur+
xHdvYP3qVcccllA8lfWjKiDUo5HuTiWMtCEmOpO6BI8mbEttroE9eBNINQxVqwZ8ZxLRqQ7m98t0
lfx0gVifCYS5LgGhOSVVU8CpywkcOr94JLM4Uvyrix4CKB5StP9QgNV3M1NrNBbTkC9Uei1ygOux
JnI/zXOMrNhQt0lsogTlXV3gSmc3NuFG87ZpeaLZETvbV5O+NamaxK4lmnujxBAzM8X4E6t0rUQT
1Y8Rcs2U5bH+nDTpTmQkq0uvz79ePD1MZjnhYffpwsXkw9e8bTdwCfRl/GEkZKdCcmPYoVO+STnB
NIJheUqThHI39AG5+MjSO7N2bpVe4pQbTNI4jqy/9/9CTLNNSWPMwoq2c92o4nBUuyRrq+QsCrlx
pPh8vkkLlGKa8cJtyV9+p5V2WMph10hXwYBlsmWDlVoqMmJB9vZPU1CRBNLXM9/yMAM1K62rhI7V
O0O3rXZBUyOiKyr+i9M1LR8vTVME+Ihrfcfr5m4YJbU9Xruc1D5zX4J/s3GkVsM8UNEe1Z2W8cDA
5VjyZ+rn3B13dg7CE8DEMUplYGYPkrfN4dIS8DwKnHKI3o/x34cKS/cyS05bveVyeJmLDwLLJqND
OKHWu0j71Q360MqkXw6+fb5QudWMiYR8Q0bjqZAU5eLjNJ0mghzuvwxw5Z5yBv4JGySyio8rAjLY
ZOXQurWTGLYijvFTOeOC3VX5hah47sYtq5zUwEMEznfm5rvv1emK5vyjYo2YtjY20tRfh8DniNoU
H7zP97iFUv/esKIpWYK+o7kF65p774du/mBjuwhKCbxUwxv1FXCSM6x21YzrbfiWk+2jD6lYa8Bz
cOMsqRIcGK5RaVPVmCSdZdvOehiE9OV3vwRAiJwGNlIzxx9lzoN/LmKgIz6dvoIxIehKeXDMHz8k
eHqHY+oPWj9V6WZBxpzp1Ti/rWICEcdL5Rmn1i62GyWfZbfNZrAPXk9MaduMT+pJ2TcvP+j6qv1g
crvB36FKNpAk7RyU9V+wupPNlF/xVGE5/D7pXUDJroq4H+qnTvnzDPCTAFqCAQWTdJ2J9nwyWRyR
hdXN3S6i+u9b1gsq405Irgd1OUyPWIp4tfFRxPPXkzGsZFGFZ+J0KLS3BszBM7y9JjCgaV9NV7M9
JyJ9eizBOYYN2jhUkcEv4SHcfSRVEy4u6y7KpM/TGM2tg9IRjiVmAa0PVSLSx90n5UptlxqF59NN
gWyf3V25BDh7Dix6O3Ax7A1rOw7tISoosnbjlJlcm9xER/xIQMch1b0vhmHYe4I4HKqo0j62QeCw
DwR+WMtq3THN6vqeA+TKU6ZjuNjg5AsyLXBvPGHs35UFhSGFa1u/U9lemOewdzJwARmhyTY3IzFc
kkv2aN+9p9DBHRtumrplFzFB+d5hQkOHz3ZaFHmzyyUtuG6UuqGmwfyJs9DL8+NVtPHlpDLQ5kqK
ypnb38WeD8IKDXIOdc+15KrmDuRb/lw045JwBtUTB7GbOfv3vPQFD4mthBbAVwqMGBexumBvxdNo
9myFucbA+jCCXMiHSmH90OqSE15OM9T7Au1IGEy15cbVgZjWfKD+1yqjG8tnmnPKegvCAIoPqKdq
yAKT0LAYCecMF5i7cENqWOaVcH4sGSEqJREaPfTwRlFvLwflPI1U7eswMkC6fPTQTko9NJBWJZM7
Ppcgxan6aZSlFzjB+KoncAth6kGXG10b/ykae1qpvzN8Q/b+vSPn3jQ/Xmbvp0iyRsJt0NJxQoTw
VqznUn51rnUrzfn2+STJr+LsuYcUKbN0rktttNNwRZym5uBBpdBcBo2zU9+lt2sH22AKBAyidsBZ
JYwjfvuhrJvgfAqxCk3eL5Dxa55+TdLSib7O0KWQbAMBLMt1PxQs0aLgXAMjZkEQgdJ/bA+6gIsQ
Qtb56RCpk3Rbqe66lWZtC6RSfZ7pwsFmG8V0xPLFgerpNupMlz4rxtV4DyLbHj42H0cTIRa3knq0
DB3dJ52Lv5EcCMlB8Th3lYLSi08diTogs69P30gVaRUB2l/PxPRspGLUsz252GKS4D00PelEm5c2
UEfv95P+TJhfRAgJ65UoC+lDFLsX90ZF9Rya7M8/HJERu3FQ9QuU3L3UdQryLXok4R4P9jq7g0BC
XqKqQ6oQJ5vS4Um13VYZ0PbWRJx0Jy4l1gRqblgdokujRFid1ihPm8Hl29T8ibRwtbbuGDp6YYHf
TNdpcbbIZGR3rBY1p3oPwSYkU4J0+5K1qfQtaf9/DenO/5fZVJImtY89Ozb/0JCPhgRn32H7xpIW
Vr5OQK06W8nmAlKURMJBJlFI1hrfYG+221b1tWY7gH+0+oA2KtZZPQCcLlz+6FukX9mzNsJEkkws
cILjKWm85xEZ2Tni3WJj9f8gdv/8YqBfjelx4tYKr9pC3cu1011nFSWxC/tyABKTDwws2jpf/05d
rQATCj2+15pVZhIJCl9csZfgAFOtCjJHhsL/DWIjKyjBivekzyU+hExLiqQBX0v1ODOp9ZV7eOQw
neNqi08O8HImsbg73/cGWjKNPJmm1JFv9sMTg6XB9qae1CM+nsVU0DpEfA6ZOWWgquFSHD1RWL9j
HD4h8VSmU/841T70AXY9ppbQLwXjw37WvdUERPA2LmcbQTZDYwxH+bUDpWlZCYi6V6NOSUdoId55
soPSye9eMchP7CZ24uDk4lQziX5O3683hhpsox99GKvwXMmFustmyfjKWYEqCwK7763h40nHiwtY
BKvE8Qmjr0QkzKwfeMTz1mlJgXHK5bc/rzOWVy9KxXXu+RlE42vY3orEhpohSamHZ4Fw9t5ISzzO
gSS25802YZBHiG1BMZhv2oiP+Weaecg2uoBEcGnUPy/DIWiZKaNlIxN4yaJHSU6+aOdswgnFr2t4
f9ael+pfPRSZ9UJbhHtNiPITYl+8Z5GfGPektraHtGVXTR6IReS38l+mMXar6QZIIhrBBeNkB5IO
FHDOtiQFpsWYtHcK8IKD2y6SQLTyXOY0hO5a9C+AwG1RpzFeva+BB4aAfhsZvK2urvxtfC6NWo3R
f7779AKYxRSIFuK0DailS/FqG/JvaJQWk9h//WuU2J/PWmVC+EdFAG6R6UNQsMWdEtL03gfWM62r
6O20G0U2CvN0JTAgQoGqkcN7OcxrokAiN++qegLrJv6B/sOx88C9KGc+vd3A8FWw2JHJUxFHy9vk
ZJnBplobhTtOxeDLkIshbEdMnA1lOBp11dCx5IuGP2L5vRde7CtvpiuJtBRCQBXQXRPUY4V34Ham
0jTQQL1eU205Yh7p0W+bvQJgj92q/CCQo83nqV88kUEVkubtoHTUpHBqI5Mdc8kBq36GL69R07L4
smmL9OvZjMsMqzqiYyUE6c3rUau3xzt0Qpv/6V2gC1HQaP0B3CEcbVztpAKDL9Im3WjWs8Fkm3Ly
QdfLrRMfAx59ccP9GYDsBLAR5RfuSOgafZZPbIpCydZLNE3j9VECZgUiHeuwKq2XXiQrMvBdZ0i+
QNCN5xuZELd27bBRuHKrvVqoRSko6io9P/3o44MqoEL+Ft02Dsz8MZIUJOH/DA4NpEynU88aTFTA
fEUsj6idlS7TgqiPKwhE/gezoR6b1r0Q8KamWzAe5f3YU7s0ewSV/f5J+sMBwD4zblyKbhxjAP8y
EhKdx53bjmlYatZGeK2yUXsmToJK0FKzZw1Kon9h19aXCML4+cm7C7rRKpCWpyonWZJoKdRbVOAz
5gmVgWmHSrVeYIH0euYN1kcS531xKem2qg+tpWiu4rb1mH012ckiRA/CBL7c4z3/2StpXALVhuWv
ttKDQBbEKoF4Ot1ThPU/UzDhPskNWHQKPITTq2GMEzuwUL6qvMubhO6jkjLJ4FfkVCrm5alw3qmz
Qgp7Ia/IoAfm8zJX+/Rsms/Cc1lwCf+m3I0q27s47FexONNXYzCO4TQ4YCNvy2LR65S9+WtkawaM
ZLh9R7J6xiwNoOdeErPt6O/tQVCBK9DtnMBCgi8cx2IMlwe/QW6GmMgJwF0gmWaCwQqNlDmn8i2l
zHTYvimgWO82wRa/uUpTjh75eP1nmGFEWjU5W3+8k77fZfNeC9qCor9+KxbwI0QWdRx5cksddfL3
Aqs4lT85PVWc90CekhRGF7ol7EY+64HC7WSO7IdGJJ7cnA4oXqmiIDTnJKBE/vdJ70kM2sLDznSF
bNhtOj4+FduSdSI81znqjOvf9vKy4sppHryVOkSzUEHQIoBmiONJBW/ZPhozrxD9CC45mjvRwflI
ilx1t7up+V2w5BZQr3GPl1d7UpXDWdC4Ku4/nrVs9qUqJq0r3oF2UAOTFUscU+2b/ZtFNT6dBtEW
LzA3dC5cnYwDiv2lnG4tKlPofc7GsXpzuH6tXlpOtXxqM7EdA663h39ry+7QhROUc1mlpK0yTwIi
wVYz17GMwSrxBfwFvOyPKe1myiZl/y/jrlbuhFoqrJJ0iFPt8FPgiJOOnJiC4YM7nd548PRVS3ge
tDTu1LY3HTy1+Y/a3seYN403PX25Uyyhl3wPbxGmTyADMHqjQrUliuQHTK5kw0xKCzr766BSgWe+
dRFGVWc+0DrRVme4dFg5CDkj2kGybN/QUsiC9kYxw/5gcU3dh12kDIlsElUPrHVezZrhwK85mun5
OIsr9+luGac8QSYCc23PIHUb0fMD9CEtc/YZAejLQ/7H8rvQerR13O5g1BS3PBxSa7uB/AKi4eBq
9ocJhZboV4UU8l2YUwDLAJ80krBLmretJBXWZ+PoJLGyRb9PRe9ez7xKg8Ik5tpQeyUgwlM7RNIi
8a1tGmC89Au9AVHsMpSeF4icvNc0fukdC5RmcYaVE4aNG07SFtpzZ1KRxfA417L32FvUWz3PNAS9
rJgreAoHKn6pzCkzgkaZ8OWDHJC3Oob7x+fRWv5jRRSL1PPXS2sjXFkGSgxVTLaYIbBdlEgshP4a
ro0i16bxT4n6jcf9zKvBGNTIZgrUseCo8rDInjUze97l6xr36RtJrtyG57iyBDmR7PZc6gVUEPzd
7TZLIiekd3Yf5CAy8S+F/52nw1tPylx6wkte8BvSdDhysOfMurZRN+/UaFql1hGUlOijJNCrbwXa
VHOCGw5y/GS5/s8K7TtGqDyl4PgsgVUqfFKywLBJxJwY4Y3btRL35HjqE/9MqVOOPx9vEtA7EXek
dNAt8n9pm9QV/wmpg2n7C7HHR3lJ31xrjG/Vbm+FPzh7I7eRV2ejpYgHtYRXBhcTZUJoDWm2euGr
t9N+4mYp1gyQy132yLOTnPfTZvclApo3PtbHBlqU+yGQz1ntThwIsGyncNWFy4tpjVlks8b71sTB
sLVgvi1bqvVJkBj+0qG0cSdFkIiM/V3xLAnybwgYxnmALaMwi9JLAFs6a6i9jHd4vFDlvwVZKOEg
ZGGnvf7j0YbP+2IcZF1/0JyufHzbprPZcmArta52K0wJWvJM44SPplOIkh/MJdqSuBdMX+p2cR6J
uWsGPwedBpOTyQtyFX/MqsO87aBOlJf+RSJa1kSFev4ph9FaQrnobozBWukPzJ+S1HkaV3dTqlCC
exfg0X40/4e7yp9+pJdtVJ+nw8ta935MlVjJG3B6JYinCmLSIoXoT4DvdGrUp6VxoQb/EU0d4hcM
KHFDxpGSR1jScxUOTexBRG/JYeoW26taTX/oO+itv/ShX6uTAGntvliiLpXpiuXmVn1lT6PGS/ur
YINDLzNDMVGVGkIx72vCi/gAkufv5MhBUO6wMUg/hejBciLEcYAWLaHSmFqYGinTxgpa8mxSaMHv
ZKAIAwVisKpY/kpBumvkStW6VbaxN7iDqR2sbEzbrg6wwjXJEK4jk8lWT1xIEEKDI51KkTMOhqzo
vIF8LGxf+Sc0J3W6/r1r6ZtZBFljr4LJfbZs0UT7sRxb2r7iQj24gbPck4tBC5o99wpoFdBEWcMZ
MBIU8UIKzlf3G3iXwtM8U3bDOgFoHqbjEQBz+Ba4WmnhyZRLHo9H6/hT7EQ6/o15dnfqjaUkp10Y
bM+kVt7cL2RhI4afR8DrADZTCVdVnxgzyyJH1TwIhD0bkGRHvP0rxmC3Tdvmm7MuswAOBLefUDm5
hiNV4/xE+QEp/f6QYl8rIWdyCuL1ftpeLCUY6wBT3zkybACEu4ShSaISXQOJVSt4t791gABH0tGL
Drt6QMQZbsGR9m7EuR+UpPuilIpUlJ6kYjNJfttFkVut1G7pQilao1d8czRtL2lXLEvgW4pzEAYJ
VQOCIxtnQoQS0164u7XyT6VX/vfZbpMxvVi9eQ1MlmhoQQ2Ne54tXFAlBTSKR3upnMt+yNvd4U8Z
StkgdCxRwyGerLh0/b0OzOiwUSdrprqkNxhrCdsQfIYLP/QwM4qaWbpqv/zRT0F3wi5FRplCiK66
ytXmm4AvPwdI2IdHVXoMhTCvnXvrKzafqWrJGSNfijsFVeP5nzCRtd67oR/0Hd+YQVcci+66MTxU
h0za5vRX//wCm0pYpoBIA2VeidohrynzIE/3XGqmvxDHgbZcJL8Yh+pnz2HP6axS5WERKaPy0PT5
ST8Dt0uyVibOVSL4eyHwniMxJDSj/mxNGJzlUBVNv/As9NaJohfrHaYEmwLbJy7LGFNTR8k/ZJDP
IffsLbjnwf7FtkovVIr2sJLV4B1xCa5twYV5tMKocpHFuofjUTpOuL1f40dvb20f+1b7OA8k+lPw
nzOxsZh+20YIVqUoLdDqyGZj8jOn/ibc9cGJoEfiZrfusd0eMMwqN3u09zbG0l+oUNzlQtHMzKdw
M9j17nW33AK8oJoTpWRyculE9twsWoJ0PBBMM1O3zlmTUXzRqsctuP1IEgkLG4S972GyrrGA4jQM
Fdm+ouv7GuBwmOgNfHmcLjt2xopC2poQunWZF5sJMTtfdIYlL+yCLq+H5XU8j5rHzKXozdV/szQU
iEB+EQ+mH1/bBBOCA4dI3JUFQWPSCfbh4sgUNpL/zGNyMhKb4fZnj9CBe3rEeffK/yat7CCHF3TK
jcjGUJuwHx1abQJ9cLy15Na19Md4WRTof7PTFZl/tZb0okcJMefd22j0TtIq+Znu8hXk/A+Hty/5
e3XThxk/dpjkLtf5yxjveSmOauSinWZgIx45nLzqlVN2x6IY9US2PdVXFXoAIBin1yYDhYrmfM4p
tIqokTNhq4b1z+fSARVl/QWUZWxhzsMPwjykuFB/3wSV+eTn6Ar+ZxKTXZ0Df+ZaYovHTDIRhfHG
eOBQCs84pQPVfxnjc/7xPpr24Db+vEA5zQrFE1bsDM19Z21OYLoIOgNRnmpmDYDZUpo3Ytdnu6gi
vomj8xQe1duLNe9iUqkzIvMwBP5jxQWthntXIl2uolmHrsdlqe7oDTD8epIPf1VDDekrofp+2Xq8
JieA3rzBCe+1I8L4pPPUZW/iH9PUYBjw+1F/gwMd1buOHNuH4LgWMi3oZONKpHb2zDn38YJTSKxQ
UaR0n5ADliRJz0VtXwIwjHiQct1LNBP7a8feWfEP+WjD2K5Y0+VEbLUfZVUUNPrtXflMIVKLxx9g
bppRM13SX85o6uqy835sGSm6w+vne24XqRRoHy7GXFFz7IkeYQwm1NdWODrImqET/vimN3Y+I9o8
dugz4tZllzv/nYHGlgE9AzhcYo/sjyyX+ce4luc84BRaV+fBNrQZWrt1LT1HvN6b5paPoIwRbpIe
yIubu4vTa9WgnNslwFOKLWM3E2ExWnOod/gPwvG5DStpNOmMULY2rPRy4uipyhXlcyRJX2tEEfSG
dHyZ8XF2esqxfRi4lPH52MYa7BJje+jBqr4s808Ox7PUUZMOwKUYETNHLkkskz6bEfAos20x4pO2
93pRnxkUNgpVyNr2q/EHcSyzZchA1UGFgYcpW4sJIhb2qUCftVDOG3XJMNgsrlyVQ75K8IAgj3hN
ttgynyEc+cnCoQ6fuZSbdXQ4FSsqtcWRgbMNdZ9+MqmfxxniKBFp2lIlptpPPveuWSv2ARJ/s9w4
WaYyzIg38ecI+U1mJ0k8+ygy0H6TlwM4tf2EM55E++w80klAs35h/lZtj2bOztoX1LlnAcRlb5AP
NNxybw2k6dtD+ZLl1Am3CD5MpIOHKtOCyKy9uGFHCcptu+CGz2bi1LeAkb2jeeMskAm+ixmyxfKs
rnLpOMi57U/vnFc1Bi3mynJlf66n6NxXFEFXOkUXozCKTVY4UB1yDWhONIEGWgeSYXZMxgSpvYkK
o79n7gY0LNtGYqZBFdaojMTjG6MzPhtFghxh0ISTgLhGRKgKrdUWuzVqNLJPK36kS1qy6xtFfyTs
QWfBT9351fhAqgWX+G3vUpmL6eKeL31eqLy64aJlV8+1iUEGbx75hcb6z7xy4sBQdhduslDB6mTB
PnezXhD9TZOLfygNOo/tcqhxhbJimsSwMFppJ1mCkVmXbB7Gtt6p+miadqhSt90a/wwx0MvXQkpR
b98ohMAVS262P5hXeJWLgHGRyBAM7t1SRYLHYNuaCYrVte8tptAxfrZYOU+df/f96F0A+fHZhP+m
2nnRnMVrWam9KO6SQg/yDdu5AJfLn6UP+E2qK+gHc132PCT/GfwXSa0oXOAu3E8KWXunegpIQwnQ
Axs66cZD5tJXRiTeZq/bbLmS27JHGvxfO+Lre9dUwC6QjPiRmXl/eHdo/HpALJLkEatC37ykmprg
OLGIdcO5e+C5+VqnZv7vH8z/4uKa+JTyJh9uC53VIypYZt9yhWy/Qq/LNTjFRIA9lOGRTqT7K+we
j7ydu0NhKKl3d1ImOBYWF7NJ7QC9BsAq18RvmWqjFNlkmaq3JZs+Bxh7vPzq/09T9jQn0VoKLzK+
xfRJBZRVUWP59l6mVSBO7Ab8Zu6SkNw1P1Vv9XnXGT4asKLahkp/W89AWQwA5k2FfhrPUuGgRkK3
C+p2nmN57mRqIN+MSBhQQftFBlg6yuIL+pnx4nHTJhPD1eMUMgnlCTiNvdnGW8hVGmzyEElgk5bS
FJebnw4NIVlBbvL3Ov9bdOR1PVnhSm24TflhFa3rbbJkzvj6wpyTh87oh8+4FCtp7R5RaPzBpJWI
p1W8Cn7qv8LbX6dAuhOYbPXnnti8omh2qzLzHAvtIObwA8sAJZ8dt8aqZY0Gct2O61qGzS09CtGx
azHld28uFe9ECDYxnAI8hMwWD5qH8cvHaQPAjrWsJFplkMybGJIk6nslsYlLwz+dsfnees3gyEEG
tQ1xAy+cRFoI5Tc5uf4kw3bgC6HmtMj9O663Q774E8FmolJFuCRcb8T3W/E0scy7j9PbmmidOJVC
4g9wFGI5ORUiF5KcK4cIPYyiBCOdFHqqPIefDuYJZzXNC3i/Re4FFTa4b56Z2oVe5dTXaivko7g+
bJezQJS19Z2Xx5BW9cJY5B6RQMgziwy5t/yEdcK/jj2CIU5AIkC7MM62hdAtg7vicqAbq9WXa2KD
i+YiV1xsxLMJ++DzRvxijv9NIC7KKOTxKltymWWR+5HeN+bLpIPvCbX1B9C4l1Ok1lFaTsZ1/XF7
N8QQQxkEzOFTb4t+caPhNga5Pj5Ir7NJ9Kh4UfEv8FaF0ayVZmIyFsiwjUuGQGSTu5GSuuv3+oVK
ZvNg/Gznjaz4vQ6kYhF7tcefZwEyBYr90RTEbsm9WT4CotQxxqaT0qW8secv8osaBHKKf8+kM2Fy
uIZu+19Vuc1BuXyRNGNAtNDNbKAmYIH1OvxbVnng0cr/GQLlaUeJinyBCHQODVss5yiz7hj+tm8S
F3hThGDG58tTf43pGa/E1pYcT2D+GdmaSdT9vc7XH8Kh0XDppB1fEPFr3ofeZ0Ml128iwLQR/6TV
u4OZNggbmiIRCYLpNfuvrujZlzvte/v3brIWYpvC7t9axwS6CJEyEFpExsvXn7GCgwUdVidxfabs
0xSkP0qA3xu2Pay5sYZqsSpz4KoOJeDY8g/0a3tc87XmdRI2TU7LQVNZp4jMk49H6T+KikFqSbp4
1aGbY4AzIywP+a5ChzbRV1twsEzH0IrS/g4LTBLou6WHkbbPy3bIaN1JQNuPB3CD4d5DwmH4IF6i
5fLb2TQJTo0zhPeGGSVM9eT0b+Uad6cR8DuA2z8/MnAjCHZwDWZaHtVjx+/c2UVgLdg8+HACQp99
9SR5KbXHtGJ0yNpRC4gTBqke6XF+Ls1JgFDgcnV5iIxTnpw28xGHMSBa6eR7YfvIhdvr1X6K9T9Z
db4c6RbcYcH5FbtHzGHEJcF6DJHZ3SOOIAgVGBVl1hu7BUe6HIMDIbcgHjTQAGlqd01rUZ49ZCZU
QZQaBANy8G5AsVQEthPyDl3Mzs8RRUd/XdLHp3Rj3BoDvLcN5TC9aBDcY8NG94Cn/HEBRGRSnVvO
zkbACmNonrP/aU7iS1WlXFym3eS1qKFyIcUChbBgNcG50qvR4tD4GLpaacDturOZbygeKlLWLSP3
LS2nT4JHhsFUlT2i+WBxRkc+uyBG59Q3Q68X6W6rGU7izNUoXCSmkyP99PHOkJPVEwVj550WoDiQ
yhsnPczG0tyMOw+e1irnHufeAAmQTIjV8tumPSTHiDjq5toWW1qf+CzP6V4NqXRE8fGBDhkt9wL+
Ah/YXXoD546zOzkNEFgHrck1ulwsGXcQG8+/POZYbsrhPzralx7GZyEKwgRqFc72HhCTp/SB7HBi
HxX8TIO04CAND8ntwTBgPiGDqydm0l8BD9A+rvwDqAqwK5C9VrpuEW7waK0pafo08ocxDrwyq98U
L2BeA6hPhtjCVj5Nl609VCLHfqkJhDFEaKqRAZiZjJaq3sZktuVYAwepkibs3Z+blCqNXsBZyAL2
7d4WsvO+IviZJi1Mg9MJ+ZjXzT5930pot/NdLdhO4ndIfUewUugeicvCi1LqgE9dUVctXZThpE87
v/K/Hbc8miMoEe2qLk7Kvl0n6oB/dK7lFewr4BwrgP+hzVdR55O3QssCrwGmHNC1yF36i6W5wxOD
4+V03O91uED+dwKwb35GDQ3wg62hQIUEEsK4LMeEvsg5Y5PtXadGWlj8VBkSRsxzQit2e1v0tiEx
I7O0i9xEAv7X/B4w5uqHAojQ7RJUkl/R80ZmJ6fniKaFEtxcvQsQskmqrVmayNITmOmoxj5o1tx8
xbPCCr/nJY5TWXzlMkWik6vZPAIjDOIKmdXg/3M/ApnkHr3tNwQm6pfHlDt+iGux5LO87quuxzLx
bQ5xVMB8aenagHLEkWvIlPZPjeQ1vn8G/4YAacxGSOKpYC010x1AwJQAU2RhhBIuU8Xitb8rFigj
shD8dZGxreWxv9JeMctT78kSu/RCJQEBlKR4XNC4fcaWYZ+K3qf71NNFIXeHFWdd2jdPx+NKzOv+
mpUzH+CufjnisGBS4fSmZ2UTEHvYUim71t89UmejTEy86TB393brNLNicLytPZeQOJ9PMefTy88s
t1lYDiPZ28NaQ7dbtUtMneaTOciQY6kZ7AZNzO3tAJ/petuJ+hjtT7tWSd60NzFDM0H/rfljkdiJ
V4VhnmNqeFSAsNby0OOqAqV2TNNqx7L3YwMz/IboO9hYyMT9AMq200uUAOQtKcfNWiAuwOqBuOlx
DW1J+O4rGy0Bbcu1sgG8U9LhtO5y1scle7HatFU2drUX9bxfFVlVtzwvcOjbCXN5a3ETagPf/EvH
V/eSFPIfFtAseQ2p+9i53MIofarAmUJ1xAzNDHibbmdij5O48UO6rqAXwLrE7xmirEV0vUqT5lW5
USJ1ILKf528zvjxbipOYssXVvkKiZDOMl5yNnu1d98/HYJlVbFbjN7fBobhSQZ3Y1bv4vhfEJX6c
Zc/s/wtcIIOKbwAdphzq4MMGHc1I+CHh5aDmc1V+x2kEjVQ88ReVZEQIgUWF9P9kocVcPSi8QmS9
kWTghO5IDO65VjNd1s5P7cccoT+tf7xOBg9yh4fq/Z41LTBfC4VHWUlYUey3GS9XxHv4BZbhvOhc
sbeKQ0yf2Go28DCQSxwaWQyRB8z6Rco7KivgWOeFROChMioBAi+5bYVGzzJdUGtqcIjDq54JiXpB
axK6ux7ryJkPtE4vgP1ZHyxK5x/fsJwH44e5KNtv4LnUhb+j7XY0QmW389Yh99Hv78YZJfbl9QfA
k6dODazzoAP2L5XkCsbz/C26Qt5c4JvbCMFyqD1Gv2T3ZfHbd+xKLv1e2Jq7BR9CZEoGv7nP/ZSW
MbnirouDvailMObGeDYYnTFJD6L4EYovNQQY18WBq/BFF87YY9R4o+hhYmu7lbNQTJkgYGiOvd91
RcIhs/AKHwFdIHHLVm9tS9e2G7HyxEi6VoFt5w/bycFutzQfPziPgjgiHBrqjXctWjNB7yI7+6Bf
cjriaqlLMnrQsBcEWCA2Chlk85HP2drpDGOsI+gVm7DtybjW9tL+cHBAhRxiOLq1o6k4VBRdbzqW
czzsWZ9/bEHPgzCW2JGxHXcGRNjlKNgvVNepLMHSxmyGx3Z19DgGcCaUKg+vjYo2n0aW9YCEo5Uq
VBdSrRykkAo1v8KsPppF7ijSZ4G505Jkzy1qZkEAIpKOYFLURdHhc87vIIi5PS197iu4fT03tCpN
zV49UG16o6ClKip2s0eIzWrqUNGzg7DzdLhVOzQuWGBGZL5nlOw6RDcvpxrudPW6FNjBCRtlotsf
2kTBC6soXVms5DTdUcJeztBQkyOh6rgQjByXZHi/UKnoz6BCLHiwHoJI00/s+UPJg8tvkw5k9+oc
QjWyR9b1aqskKP7ez41jhKNwWRfkeFS/fsGnG9a8BMhdQ/NStZtKt9QRbdoe1hVHWcE1H0CaZNxQ
T2HFqM9XNoUtiegbjtXoVhX6K6mfI6z163eR6NyEuNgDFQTJcLbmZLfFnNTqe9UQSHr7Y452nrn5
4+1t0/sPgkUBxncXuJmM/Ud9nsB5gOI2GOic2KOE+Am7ns1nTrqimTA9e1ZnspbxakpPT0KEhAcC
0I6LpYk8DxyH2+Fn5pTASDDedsTIl89HECzGd0VA1b3ccFCckb3ylRi2lXzD7qf43UN9ctoEtlJ9
FGpVieIMavexgcH8qn42oECi+WZkosXJWCmxdIkD1PYVhtn+8jLzPMzlbXCdPUserrtt6tPlrG9e
lEfj+MSl6KVki7pXJIYPMPca+uJoJrJF13BLcAC1eu9hG/mSy/9r7SHJ4mhb/lES1nUI5RwzIp+i
wtJ8NmWu905idTy9mA4jN5tuI3m3cRTskLrQYFMHPw6ORhIzbq7zXqpMDxb2tvzTOW1CE5I+KuUH
CcV/TA9ccX3miwi5XlYk8hMq6lWxJuRScrBf/ldixaHWmgHRBLEWQod4TBJFl4lPhCSTOiWH0mQp
jKAKKGue4nPknUKJXYg1dteDSZ02/d+F69c8XWyRJymD5UuORmXgeN+LOalBwIrNHrdJgPbCnx4y
IoJt9WK+Xo0Bmmra1jn7U1wP7DnqCAqs/HQ6INQS9cyoMU5NC5V8ndAZvYNPKsTItLNAgUDjSKHy
+WJzqTUc9hpFZUawj2PDq+kqPcvK/xF3cpIEmYMsF63f9iOyN0ignAIPPcyOjXiYPn5/Ap6dXD0Y
jtrtV8EBGMDiIatDJlJ7nzuKSgZeF1QTDZKfqJkDrc3SldIehuBvYbe0kvXUUOhVYZqynm4u+UrV
b0E3O+HWcclcQafxMdII60ykBg3PSAeOJO8C74VzF2guZISUPE4CxkWMI1sEDGGrxjGuV13bWac5
a+/nQaxBzY3SokHXYGxkw8MFKH14TV119621O0R+e7Y4ehEI8C+47nd36z7iPObO9tZS16dVKf2X
sDSzQEdpRTg/OUEPOFvO0ncXq1oT4QpXyC/exUoYg8tCvLKd/Gyzyz5KVlzvokdv7QTTrFgU+cb+
LUKwORrGm71+v+J9p8YwfuFQkCCCl3A1tc/EMBzvc3RUEdZoRPo6IKbnePVx6oeQUEOZD7CTr0YV
Jo84KeUEIEQ0jaCrkxOBs2EuZsST2QOxpoV/VwCLInW9MI7Iv15i/bRq5fLN6Ip61C33IRAQ70j1
u9VjkXbjoZsYmfQMRjof8iXBMZjKQQ0MHhFOSyDMWRj7PjfXwcxEMRo/h4fnj3JHksq+nCZs53y+
4KPdQXPr6iJkDPEQpNKr9GkrlQKr4paxj2fFxusiTDQCHYczqa8/u8NjnAlBxGdqaDTt+LDKaLIb
O8z630zP/pHHM7KB4fH220lfFQRILvtFN83b+tGoo3cs+fmVeA+7joQW5WFKENeZ++Bysg91ovh0
F70iqiyhNC23nQpSWdwzGZMnmHi3sspih/+ECQmmPVfRwURrpRg9JycS+Z+d1dFLSN+SAmFpq/U/
/i0iAk2ljG3FjSACbRiN6L0IEvuN3PeUKucd32qTSChJyWZlv8VTND5zEdHRu8Cu+UgOu3jUqQEp
cnPkUPrVTdrnhem4mRL+MlfvB/c8xDUWAtcUyg1z7njUL/0DHW8TBfgBlLbT0SNXekQzPuZyF9BW
kzY3Wku3a9p/OuiPhCNGTCBbl/xurPdiuQrxxeX+0GXBgxH9LFG2Vjlz4SnZhU0QZ8sIigFFlmt2
vw80Z8BpDpXrmXVLUVMH2zB1qZVm9KxZHLJc//nWg0UJBIyyTkwgg0hginLdWa/jiIg23C7zkpkG
pf/QK+r0xb66MSC7/QSrXGH6zKwUO3swT4k96cZsECCzmzRtT3jIYGkUXRVfacAFoGIzqOExIlDw
PfLKyFoSqcDT7nxT+h4f6aJPIGxvr219cNsEdrTjw92h2YugLkphD130zUS6LTefbCEWXsenks2g
VsZzUm9aFSLSh6W9GXr40hY0MWle2WM1onADc4jDYyzEfpSx7Ny78z00ogOi5pQyXBcbno5hykAU
V1qTnlbEh4jwMU/OJFk+F8cvOp0h9lGlhOe+CUQzaLYE9LnIwTknXOFvReVfraw7whIwLCi2P618
S/40Z5cqf3vkmejN9jbD6HICSam4MHRJzw==
`protect end_protected
